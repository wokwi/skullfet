magic
tech sky130A
timestamp 1699107033
<< obsm1 >>
rect 0 950 7850 2550
<< obsm2 >>
rect 0 950 7850 2550
<< obsm3 >>
rect 0 950 7850 2550
<< obsm4 >>
rect 0 950 7850 2550
<< metal3 >>
rect 0 0 2400 150
rect 5450 0 7850 150
<< metal4 >>
rect 520 2330 1160 2410
rect 1560 2330 1640 2410
rect 1960 2330 2040 2410
rect 440 2250 1160 2330
rect 1480 2250 1640 2330
rect 1880 2250 2120 2330
rect 360 1770 600 2250
rect 920 2090 1160 2250
rect 920 2010 1080 2090
rect 920 1930 1000 2010
rect 1400 1930 1640 2250
rect 1800 2170 2120 2250
rect 1720 2090 2040 2170
rect 1720 2010 1960 2090
rect 1720 1930 1880 2010
rect 1400 1850 1880 1930
rect 1320 1770 1800 1850
rect 200 1690 1160 1770
rect 1240 1690 1800 1770
rect 280 1610 1160 1690
rect 520 1370 600 1450
rect 440 1290 600 1370
rect 920 1290 1160 1610
rect 1400 1610 1880 1690
rect 360 1210 1080 1290
rect 280 1130 1000 1210
rect 1400 1130 1640 1610
rect 1720 1530 1880 1610
rect 1720 1450 1960 1530
rect 1720 1370 2040 1450
rect 1800 1290 2120 1370
rect 1880 1210 2120 1290
rect 2200 1290 2440 2410
rect 2760 2330 2840 2410
rect 3240 2330 3320 2410
rect 4040 2330 4120 2410
rect 5000 2330 5640 2410
rect 6040 2330 6680 2410
rect 2760 2250 2920 2330
rect 3160 2250 3320 2330
rect 3960 2250 4120 2330
rect 4920 2250 5640 2330
rect 5960 2250 6680 2330
rect 7080 2250 7320 2410
rect 2760 1290 3000 2250
rect 3080 1290 3320 2250
rect 3720 1290 3800 1370
rect 2200 1210 2920 1290
rect 3080 1210 3480 1290
rect 3640 1210 3800 1290
rect 1960 1130 2040 1210
rect 2200 1130 2840 1210
rect 3080 1130 3800 1210
rect 3880 1290 4120 2250
rect 4840 1850 5080 2250
rect 5400 2090 5640 2250
rect 5400 2010 5560 2090
rect 5400 1930 5480 2010
rect 5880 1850 6120 2250
rect 6440 2090 6680 2250
rect 6760 2170 7560 2250
rect 6840 2090 7640 2170
rect 6440 2010 6600 2090
rect 7000 2010 7640 2090
rect 6440 1930 6520 2010
rect 4760 1770 5320 1850
rect 5800 1770 6360 1850
rect 4680 1690 5320 1770
rect 5720 1690 6360 1770
rect 4520 1290 4600 1370
rect 3880 1210 4280 1290
rect 4440 1210 4600 1290
rect 3880 1130 4600 1210
rect 4840 1130 5080 1690
rect 5880 1290 6120 1690
rect 6440 1530 6520 1610
rect 6440 1450 6600 1530
rect 6440 1290 6680 1450
rect 5880 1130 6680 1290
rect 7080 1290 7320 2010
rect 7480 1930 7640 2010
rect 7560 1850 7640 1930
rect 7080 1210 7480 1290
rect 7000 1130 7400 1210
rect 1400 1050 1480 1130
rect 3080 1050 3160 1130
rect 3880 1050 3960 1130
<< labels >>
flabel metal3 s 0 0 2400 150 0 FreeSans 240 0 0 0 VPWR
port 1 nsew power input
flabel metal3 s 5450 0 7850 150 0 FreeSans 240 0 0 0 VGND
port 2 nsew ground input
<< end >>
