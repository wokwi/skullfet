magic
tech sky130A
timestamp 1638034600
<< metal1 >>
rect 30 -20 40 -10
rect 40 -20 50 0
rect 50 -20 60 0
rect 60 -20 70 0
rect 70 -20 80 0
rect 80 -20 90 0
rect 90 -20 100 0
rect 100 -20 110 0
rect 110 -20 120 0
rect 160 -20 170 -10
rect 170 -20 180 0
rect 210 -20 220 -10
rect 220 -20 230 0
rect 230 -20 240 -10
rect 250 -20 260 0
rect 260 -20 270 0
rect 270 -20 280 0
rect 320 -20 330 0
rect 330 -20 340 -10
rect 370 -20 380 -10
rect 380 -20 390 0
rect 470 -20 480 -10
rect 480 -20 490 0
rect 590 -20 600 -10
rect 600 -20 610 0
rect 610 -20 620 0
rect 620 -20 630 0
rect 630 -20 640 0
rect 640 -20 650 0
rect 650 -20 660 0
rect 660 -20 670 0
rect 670 -20 680 0
rect 720 -20 730 -10
rect 730 -20 740 0
rect 740 -20 750 0
rect 750 -20 760 0
rect 760 -20 770 0
rect 770 -20 780 0
rect 780 -20 790 0
rect 790 -20 800 0
rect 800 -20 810 0
rect 860 -20 870 0
rect 870 -20 880 0
rect 880 -20 890 0
rect 20 -40 30 -20
rect 30 -40 40 -20
rect 40 -40 50 -20
rect 90 -40 100 -20
rect 100 -40 110 -20
rect 110 -40 120 -20
rect 150 -40 160 -20
rect 160 -40 170 -20
rect 170 -40 180 -20
rect 190 -40 200 -30
rect 200 -40 210 -20
rect 210 -40 220 -20
rect 220 -40 230 -20
rect 230 -30 240 -20
rect 250 -40 260 -20
rect 260 -40 270 -20
rect 270 -40 280 -20
rect 320 -40 330 -20
rect 330 -40 340 -20
rect 340 -40 350 -20
rect 360 -40 370 -20
rect 370 -40 380 -20
rect 380 -40 390 -20
rect 460 -40 470 -20
rect 470 -40 480 -20
rect 480 -40 490 -20
rect 580 -40 590 -20
rect 590 -40 600 -20
rect 600 -40 610 -20
rect 650 -40 660 -20
rect 660 -40 670 -20
rect 670 -40 680 -20
rect 710 -40 720 -20
rect 720 -40 730 -20
rect 730 -40 740 -20
rect 780 -40 790 -20
rect 790 -40 800 -20
rect 800 -40 810 -20
rect 820 -30 830 -20
rect 830 -40 840 -20
rect 840 -40 850 -20
rect 850 -40 860 -20
rect 860 -40 870 -20
rect 870 -40 880 -20
rect 880 -40 890 -20
rect 890 -40 900 -20
rect 900 -40 910 -20
rect 910 -40 920 -20
rect 920 -40 930 -30
rect 20 -60 30 -40
rect 30 -60 40 -40
rect 40 -60 50 -40
rect 90 -60 100 -40
rect 100 -50 110 -40
rect 150 -60 160 -40
rect 160 -60 170 -40
rect 170 -60 180 -40
rect 190 -60 200 -40
rect 200 -60 210 -40
rect 210 -50 220 -40
rect 250 -60 260 -40
rect 260 -60 270 -40
rect 270 -60 280 -40
rect 320 -60 330 -40
rect 330 -60 340 -40
rect 340 -60 350 -40
rect 360 -60 370 -40
rect 370 -60 380 -40
rect 380 -60 390 -40
rect 460 -60 470 -40
rect 470 -60 480 -40
rect 480 -60 490 -40
rect 580 -60 590 -40
rect 590 -60 600 -40
rect 600 -60 610 -40
rect 650 -60 660 -40
rect 660 -50 670 -40
rect 710 -60 720 -40
rect 720 -60 730 -40
rect 730 -60 740 -40
rect 780 -60 790 -40
rect 790 -50 800 -40
rect 850 -50 860 -40
rect 860 -60 870 -40
rect 870 -60 880 -40
rect 880 -60 890 -40
rect 890 -50 900 -40
rect 900 -50 910 -40
rect 910 -60 920 -40
rect 920 -60 930 -40
rect 20 -80 30 -60
rect 30 -80 40 -60
rect 40 -80 50 -60
rect 140 -80 150 -70
rect 150 -80 160 -60
rect 160 -80 170 -60
rect 170 -80 180 -60
rect 180 -80 190 -60
rect 190 -80 200 -60
rect 200 -70 210 -60
rect 250 -80 260 -60
rect 260 -80 270 -60
rect 270 -80 280 -60
rect 320 -80 330 -60
rect 330 -80 340 -60
rect 340 -80 350 -60
rect 360 -80 370 -60
rect 370 -80 380 -60
rect 380 -80 390 -60
rect 460 -80 470 -60
rect 470 -80 480 -60
rect 480 -80 490 -60
rect 570 -80 580 -70
rect 580 -80 590 -60
rect 590 -80 600 -60
rect 600 -80 610 -60
rect 610 -80 620 -70
rect 620 -80 630 -70
rect 630 -80 640 -70
rect 700 -80 710 -70
rect 710 -80 720 -60
rect 720 -80 730 -60
rect 730 -80 740 -60
rect 740 -80 750 -70
rect 750 -80 760 -70
rect 760 -80 770 -70
rect 860 -80 870 -60
rect 870 -80 880 -60
rect 880 -80 890 -60
rect 920 -70 930 -60
rect 0 -90 10 -80
rect 10 -100 20 -80
rect 20 -100 30 -80
rect 30 -100 40 -80
rect 40 -100 50 -80
rect 50 -100 60 -80
rect 60 -100 70 -80
rect 70 -100 80 -80
rect 80 -100 90 -80
rect 90 -100 100 -80
rect 100 -100 110 -80
rect 110 -100 120 -80
rect 130 -90 140 -80
rect 140 -90 150 -80
rect 150 -100 160 -80
rect 160 -100 170 -80
rect 170 -100 180 -80
rect 180 -100 190 -80
rect 190 -100 200 -80
rect 200 -100 210 -90
rect 250 -100 260 -80
rect 260 -100 270 -80
rect 270 -100 280 -80
rect 320 -100 330 -80
rect 330 -100 340 -80
rect 340 -100 350 -80
rect 360 -100 370 -80
rect 370 -100 380 -80
rect 380 -100 390 -80
rect 460 -100 470 -80
rect 470 -100 480 -80
rect 480 -100 490 -80
rect 560 -90 570 -80
rect 570 -90 580 -80
rect 580 -100 590 -80
rect 590 -100 600 -80
rect 600 -100 610 -80
rect 610 -90 620 -80
rect 620 -90 630 -80
rect 630 -90 640 -80
rect 690 -90 700 -80
rect 700 -90 710 -80
rect 710 -100 720 -80
rect 720 -100 730 -80
rect 730 -100 740 -80
rect 740 -90 750 -80
rect 750 -90 760 -80
rect 760 -90 770 -80
rect 860 -100 870 -80
rect 870 -100 880 -80
rect 880 -100 890 -80
rect 90 -120 100 -100
rect 100 -120 110 -100
rect 110 -120 120 -100
rect 150 -120 160 -100
rect 160 -120 170 -100
rect 170 -120 180 -100
rect 190 -120 200 -100
rect 200 -120 210 -100
rect 210 -120 220 -110
rect 250 -120 260 -100
rect 260 -120 270 -100
rect 270 -120 280 -100
rect 320 -120 330 -100
rect 330 -120 340 -100
rect 340 -120 350 -100
rect 360 -120 370 -100
rect 370 -120 380 -100
rect 380 -120 390 -100
rect 460 -120 470 -100
rect 470 -120 480 -100
rect 480 -120 490 -100
rect 580 -120 590 -100
rect 590 -120 600 -100
rect 600 -120 610 -100
rect 710 -120 720 -100
rect 720 -120 730 -100
rect 730 -120 740 -100
rect 780 -120 790 -100
rect 790 -120 800 -110
rect 860 -120 870 -100
rect 870 -120 880 -100
rect 880 -120 890 -100
rect 30 -140 40 -130
rect 40 -140 50 -120
rect 90 -140 100 -120
rect 100 -140 110 -120
rect 110 -140 120 -120
rect 150 -140 160 -120
rect 160 -140 170 -120
rect 170 -140 180 -120
rect 190 -130 200 -120
rect 200 -140 210 -120
rect 210 -140 220 -120
rect 220 -140 230 -120
rect 230 -140 240 -130
rect 250 -140 260 -120
rect 260 -140 270 -120
rect 270 -140 280 -120
rect 320 -140 330 -120
rect 330 -140 340 -120
rect 340 -140 350 -120
rect 360 -140 370 -120
rect 370 -140 380 -120
rect 380 -140 390 -120
rect 440 -140 450 -130
rect 460 -140 470 -120
rect 470 -140 480 -120
rect 480 -140 490 -120
rect 540 -140 550 -130
rect 580 -140 590 -120
rect 590 -140 600 -120
rect 600 -140 610 -120
rect 710 -140 720 -120
rect 720 -140 730 -120
rect 730 -140 740 -120
rect 780 -140 790 -120
rect 790 -140 800 -120
rect 800 -140 810 -120
rect 860 -140 870 -120
rect 870 -140 880 -120
rect 880 -140 890 -120
rect 10 -160 20 -150
rect 20 -160 30 -140
rect 30 -160 40 -140
rect 40 -160 50 -140
rect 50 -160 60 -140
rect 60 -160 70 -140
rect 70 -160 80 -140
rect 80 -160 90 -140
rect 90 -160 100 -140
rect 100 -150 110 -140
rect 150 -160 160 -140
rect 160 -160 170 -140
rect 170 -160 180 -140
rect 210 -150 220 -140
rect 220 -160 230 -140
rect 230 -150 240 -140
rect 250 -160 260 -140
rect 260 -160 270 -140
rect 270 -160 280 -140
rect 280 -160 290 -140
rect 290 -160 300 -140
rect 300 -160 310 -140
rect 310 -160 320 -140
rect 320 -160 330 -140
rect 330 -150 340 -140
rect 360 -160 370 -140
rect 370 -160 380 -140
rect 380 -160 390 -140
rect 390 -160 400 -140
rect 400 -160 410 -140
rect 410 -160 420 -150
rect 420 -160 430 -150
rect 430 -160 440 -140
rect 440 -160 450 -140
rect 460 -160 470 -140
rect 470 -160 480 -140
rect 480 -160 490 -140
rect 490 -160 500 -140
rect 500 -160 510 -140
rect 510 -160 520 -150
rect 520 -160 530 -150
rect 530 -160 540 -140
rect 540 -160 550 -140
rect 580 -160 590 -140
rect 590 -160 600 -140
rect 600 -160 610 -140
rect 710 -160 720 -140
rect 720 -160 730 -140
rect 730 -160 740 -140
rect 740 -160 750 -140
rect 750 -160 760 -140
rect 760 -160 770 -140
rect 770 -160 780 -140
rect 780 -160 790 -140
rect 790 -160 800 -140
rect 800 -160 810 -140
rect 850 -160 860 -150
rect 860 -160 870 -140
rect 870 -160 880 -140
rect 880 -160 890 -140
rect 890 -160 900 -140
rect 900 -150 910 -140
rect 150 -170 160 -160
rect 360 -170 370 -160
rect 460 -170 470 -160
<< end >>
