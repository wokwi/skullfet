magic
tech sky130A
magscale 1 2
timestamp 1640767452
<< nwell >>
rect 2187 1269 3240 2025
rect 1134 1053 3240 1269
rect 1134 216 2106 1053
<< nmos >>
rect 1215 2403 2025 2511
rect 351 1161 459 1971
<< pmos >>
rect 2781 1161 2889 1971
rect 1215 567 2025 675
<< ndiff >>
rect 1431 2727 1863 2781
rect 1377 2673 1863 2727
rect 1269 2646 1971 2673
rect 1269 2592 1296 2646
rect 1350 2592 1971 2646
rect 1269 2565 1971 2592
rect 1215 2511 2025 2565
rect 1215 2349 2025 2403
rect 1215 2295 1377 2349
rect 1215 2241 1323 2295
rect 1269 2187 1323 2241
rect 1539 2187 1701 2349
rect 1863 2295 1944 2349
rect 1998 2295 2025 2349
rect 1917 2241 2025 2295
rect 1917 2187 1971 2241
rect 1269 2133 1377 2187
rect 1485 2133 1755 2187
rect 1863 2133 1971 2187
rect 1269 2079 1593 2133
rect 1647 2079 1917 2133
rect 1377 2025 1539 2079
rect 1701 2025 1917 2079
rect 297 1917 351 1971
rect 189 1809 351 1917
rect 81 1377 351 1809
rect 135 1323 351 1377
rect 189 1296 351 1323
rect 189 1242 216 1296
rect 270 1242 351 1296
rect 189 1215 351 1242
rect 297 1161 351 1215
rect 459 1944 621 1971
rect 459 1890 513 1944
rect 567 1917 621 1944
rect 1431 1917 1809 2025
rect 567 1890 729 1917
rect 459 1863 729 1890
rect 1431 1863 1485 1917
rect 1539 1863 1593 1917
rect 1647 1863 1701 1917
rect 1755 1863 1809 1917
rect 459 1809 567 1863
rect 675 1809 837 1863
rect 459 1647 513 1809
rect 729 1755 837 1809
rect 729 1701 999 1755
rect 675 1647 945 1701
rect 459 1593 783 1647
rect 837 1593 999 1647
rect 459 1539 729 1593
rect 837 1539 945 1593
rect 459 1485 783 1539
rect 837 1485 999 1539
rect 459 1323 513 1485
rect 675 1431 945 1485
rect 729 1377 999 1431
rect 729 1323 837 1377
rect 459 1269 567 1323
rect 675 1269 783 1323
rect 459 1215 783 1269
rect 459 1161 621 1215
<< pdiff >>
rect 2619 1944 2781 1971
rect 2619 1917 2673 1944
rect 2457 1890 2673 1917
rect 2727 1890 2781 1944
rect 2457 1863 2781 1890
rect 2457 1809 2565 1863
rect 2673 1809 2781 1863
rect 2403 1755 2511 1809
rect 2241 1701 2511 1755
rect 2295 1647 2565 1701
rect 2727 1647 2781 1809
rect 2241 1593 2403 1647
rect 2457 1593 2781 1647
rect 2295 1539 2403 1593
rect 2511 1539 2781 1593
rect 2241 1485 2403 1539
rect 2457 1485 2781 1539
rect 2295 1431 2565 1485
rect 2241 1377 2511 1431
rect 2403 1323 2511 1377
rect 2727 1323 2781 1485
rect 2403 1269 2565 1323
rect 2673 1269 2781 1323
rect 2511 1242 2781 1269
rect 2511 1215 2673 1242
rect 1431 1161 1485 1215
rect 1539 1161 1593 1215
rect 1647 1161 1701 1215
rect 1755 1161 1809 1215
rect 2619 1188 2673 1215
rect 2727 1188 2781 1242
rect 2619 1161 2781 1188
rect 2889 1917 2943 1971
rect 2889 1809 3051 1917
rect 2889 1755 3105 1809
rect 2889 1323 3159 1755
rect 2889 1296 3051 1323
rect 2889 1242 2970 1296
rect 3024 1242 3051 1296
rect 2889 1215 3051 1242
rect 2889 1161 2943 1215
rect 1431 1053 1809 1161
rect 1377 999 1539 1053
rect 1701 999 1917 1053
rect 1269 945 1593 999
rect 1647 945 1917 999
rect 1269 891 1377 945
rect 1485 891 1755 945
rect 1863 891 1971 945
rect 1269 837 1323 891
rect 1215 783 1323 837
rect 1215 729 1377 783
rect 1539 729 1701 891
rect 1917 837 1971 891
rect 1917 783 2025 837
rect 1863 729 1944 783
rect 1998 729 2025 783
rect 1215 675 2025 729
rect 1215 513 2025 567
rect 1269 486 1971 513
rect 1269 432 1890 486
rect 1944 432 1971 486
rect 1269 405 1971 432
rect 1377 351 1863 405
rect 1431 297 1863 351
<< ndiffc >>
rect 1296 2592 1350 2646
rect 1944 2295 1998 2349
rect 216 1242 270 1296
rect 513 1890 567 1944
<< pdiffc >>
rect 2673 1890 2727 1944
rect 2673 1188 2727 1242
rect 2970 1242 3024 1296
rect 1944 729 1998 783
rect 1890 432 1944 486
<< psubdiff >>
rect 27 1242 135 1269
rect 27 1161 81 1242
rect 27 1134 135 1161
<< nsubdiff >>
rect 3105 1242 3186 1269
rect 3159 1161 3186 1242
rect 3105 1107 3186 1161
rect 1917 297 1944 351
rect 2025 297 2052 351
rect 1917 270 2052 297
<< psubdiffcont >>
rect 81 1161 135 1242
<< nsubdiffcont >>
rect 3105 1161 3159 1242
rect 1944 297 2025 351
<< poly >>
rect 1053 2403 1215 2511
rect 2025 2484 2889 2511
rect 2025 2430 2376 2484
rect 2430 2430 2808 2484
rect 2862 2430 2889 2484
rect 2025 2403 2889 2430
rect 351 1971 459 2133
rect 2781 1971 2889 2403
rect 351 675 459 1161
rect 2781 999 2889 1161
rect 351 648 1215 675
rect 351 594 378 648
rect 432 594 810 648
rect 864 594 1215 648
rect 351 567 1215 594
rect 2025 567 2187 675
<< polycont >>
rect 2376 2430 2430 2484
rect 2808 2430 2862 2484
rect 378 594 432 648
rect 810 594 864 648
<< locali >>
rect 486 2646 1350 2673
rect 486 2592 1296 2646
rect 486 2565 1350 2592
rect 486 1944 594 2565
rect 2349 2484 2889 2511
rect 2349 2430 2376 2484
rect 2430 2430 2808 2484
rect 2862 2430 2889 2484
rect 2349 2403 2889 2430
rect 1944 2349 2295 2376
rect 1998 2295 2295 2349
rect 1944 2268 2295 2295
rect 2187 2160 2754 2268
rect 486 1890 513 1944
rect 567 1890 594 1944
rect 2646 1944 2754 2160
rect 2646 1890 2673 1944
rect 2727 1890 2754 1944
rect 81 1242 216 1296
rect 270 1242 297 1296
rect 2943 1242 2970 1296
rect 3024 1269 3051 1296
rect 3024 1242 3159 1269
rect 135 1161 297 1242
rect 81 1134 297 1161
rect 189 513 297 1134
rect 2646 1188 2673 1242
rect 2727 1188 2754 1242
rect 2646 810 2754 1188
rect 1944 783 2754 810
rect 1998 729 2754 783
rect 1944 702 2754 729
rect 2943 1161 3105 1242
rect 2943 1134 3159 1161
rect 351 648 891 675
rect 351 594 378 648
rect 432 594 810 648
rect 864 594 891 648
rect 351 567 891 594
rect 2943 594 3051 1134
rect 189 405 216 513
rect 1890 486 2349 513
rect 1944 432 2349 486
rect 1890 405 2349 432
rect 2430 405 3051 513
rect 1890 351 2079 405
rect 1890 297 1944 351
rect 2025 297 2079 351
<< viali >>
rect 2943 513 3051 594
rect 216 405 297 513
rect 2349 405 2430 513
<< metal1 >>
rect 1431 2727 1863 2781
rect 1377 2673 1863 2727
rect 1269 2565 1971 2673
rect 1215 2349 2025 2565
rect 1215 2295 1377 2349
rect 1215 2241 1323 2295
rect 1269 2187 1323 2241
rect 1539 2187 1701 2349
rect 1863 2295 2025 2349
rect 1917 2241 2025 2295
rect 1917 2187 1971 2241
rect 1269 2133 1377 2187
rect 1485 2133 1755 2187
rect 1863 2133 1971 2187
rect 1269 2079 1593 2133
rect 1647 2079 1917 2133
rect 1377 2025 1539 2079
rect 1701 2025 1917 2079
rect 297 1917 621 1971
rect 1431 1917 1809 2025
rect 2619 1917 2943 1971
rect 189 1863 729 1917
rect 1107 1863 1269 1917
rect 1431 1863 1485 1917
rect 1539 1863 1593 1917
rect 1647 1863 1701 1917
rect 1755 1863 1809 1917
rect 1971 1863 2133 1917
rect 2457 1863 3051 1917
rect 189 1809 567 1863
rect 675 1809 837 1863
rect 81 1647 513 1809
rect 729 1755 837 1809
rect 1053 1755 1323 1863
rect 1917 1755 2187 1863
rect 2457 1809 2565 1863
rect 2673 1809 3051 1863
rect 2403 1755 2511 1809
rect 729 1701 999 1755
rect 1107 1701 1431 1755
rect 1809 1701 2133 1755
rect 2241 1701 2511 1755
rect 2727 1755 3105 1809
rect 675 1647 945 1701
rect 1269 1647 1485 1701
rect 1755 1647 1971 1701
rect 2295 1647 2565 1701
rect 2727 1647 3159 1755
rect 81 1593 783 1647
rect 837 1593 999 1647
rect 1377 1593 1593 1647
rect 1647 1593 1863 1647
rect 2241 1593 2403 1647
rect 2457 1593 3159 1647
rect 81 1539 729 1593
rect 837 1539 945 1593
rect 81 1485 783 1539
rect 837 1485 999 1539
rect 1485 1485 1755 1593
rect 2295 1539 2403 1593
rect 2511 1539 3159 1593
rect 2241 1485 2403 1539
rect 2457 1485 3159 1539
rect 81 1377 513 1485
rect 675 1431 945 1485
rect 1377 1431 1593 1485
rect 1647 1431 1863 1485
rect 2295 1431 2565 1485
rect 135 1323 513 1377
rect 729 1377 999 1431
rect 1107 1377 1485 1431
rect 1755 1377 2187 1431
rect 2241 1377 2511 1431
rect 729 1323 837 1377
rect 1053 1323 1377 1377
rect 1863 1323 2187 1377
rect 189 1269 567 1323
rect 675 1269 783 1323
rect 189 1215 783 1269
rect 1053 1269 1269 1323
rect 1971 1269 2187 1323
rect 2403 1323 2511 1377
rect 2727 1323 3159 1485
rect 2403 1269 2565 1323
rect 2673 1269 3051 1323
rect 1053 1215 1215 1269
rect 2025 1215 2187 1269
rect 2511 1215 3051 1269
rect 297 1161 621 1215
rect 1107 1161 1161 1215
rect 1431 1161 1485 1215
rect 1539 1161 1593 1215
rect 1647 1161 1701 1215
rect 1755 1161 1809 1215
rect 2079 1161 2133 1215
rect 2619 1161 2943 1215
rect 1431 1053 1809 1161
rect 1377 999 1539 1053
rect 1701 999 1917 1053
rect 1269 945 1593 999
rect 1647 945 1917 999
rect 1269 891 1377 945
rect 1485 891 1755 945
rect 1863 891 1971 945
rect 1269 837 1323 891
rect 1215 783 1323 837
rect 1215 729 1377 783
rect 1539 729 1701 891
rect 1917 837 1971 891
rect 1917 783 2025 837
rect 1863 729 2025 783
rect 189 513 621 540
rect 1215 513 2025 729
rect 2322 594 3132 621
rect 2322 513 2943 594
rect 3051 513 3132 594
rect 189 405 216 513
rect 297 405 621 513
rect 1269 405 1971 513
rect 2322 405 2349 513
rect 2430 405 3132 513
rect 189 378 621 405
rect 189 216 297 378
rect 1377 351 1863 405
rect 2322 351 3132 405
rect 1431 297 1863 351
rect 0 135 2943 216
rect 3024 81 3132 351
rect 0 0 3132 81
<< metal2 >>
rect 1431 2727 1863 2781
rect 1377 2673 1863 2727
rect 1269 2565 1971 2673
rect 1215 2349 2025 2565
rect 1215 2295 1377 2349
rect 1215 2241 1323 2295
rect 1269 2187 1323 2241
rect 1539 2187 1701 2349
rect 1863 2295 2025 2349
rect 1917 2241 2025 2295
rect 1917 2187 1971 2241
rect 1269 2133 1377 2187
rect 1485 2133 1755 2187
rect 1863 2133 1971 2187
rect 1269 2079 1593 2133
rect 1647 2079 1917 2133
rect 1377 2025 1539 2079
rect 1701 2025 1917 2079
rect 297 1917 621 1971
rect 1431 1917 1809 2025
rect 2619 1917 2943 1971
rect 189 1863 729 1917
rect 1431 1863 1485 1917
rect 1539 1863 1593 1917
rect 1647 1863 1701 1917
rect 1755 1863 1809 1917
rect 2457 1863 3051 1917
rect 189 1809 567 1863
rect 675 1809 837 1863
rect 2457 1809 2565 1863
rect 2673 1809 3051 1863
rect 81 1647 513 1809
rect 729 1755 837 1809
rect 2403 1755 2511 1809
rect 729 1701 999 1755
rect 2241 1701 2511 1755
rect 2727 1755 3105 1809
rect 675 1647 945 1701
rect 2295 1647 2565 1701
rect 2727 1647 3159 1755
rect 81 1593 783 1647
rect 837 1593 999 1647
rect 2241 1593 2403 1647
rect 2457 1593 3159 1647
rect 81 1539 729 1593
rect 837 1539 945 1593
rect 2295 1539 2403 1593
rect 2511 1539 3159 1593
rect 81 1485 783 1539
rect 837 1485 999 1539
rect 2241 1485 2403 1539
rect 2457 1485 3159 1539
rect 81 1377 513 1485
rect 675 1431 945 1485
rect 2295 1431 2565 1485
rect 135 1323 513 1377
rect 729 1377 999 1431
rect 2241 1377 2511 1431
rect 729 1323 837 1377
rect 2403 1323 2511 1377
rect 2727 1323 3159 1485
rect 189 1269 567 1323
rect 675 1269 783 1323
rect 2403 1269 2565 1323
rect 2673 1269 3051 1323
rect 189 1215 783 1269
rect 2511 1215 3051 1269
rect 297 1161 621 1215
rect 1431 1161 1485 1215
rect 1539 1161 1593 1215
rect 1647 1161 1701 1215
rect 1755 1161 1809 1215
rect 2619 1161 2943 1215
rect 1431 1053 1809 1161
rect 1377 999 1539 1053
rect 1701 999 1917 1053
rect 1269 945 1593 999
rect 1647 945 1917 999
rect 1269 891 1377 945
rect 1485 891 1755 945
rect 1863 891 1971 945
rect 1269 837 1323 891
rect 1215 783 1323 837
rect 1215 729 1377 783
rect 1539 729 1701 891
rect 1917 837 1971 891
rect 1917 783 2025 837
rect 1863 729 2025 783
rect 1215 513 2025 729
rect 1269 405 1971 513
rect 1377 351 1863 405
rect 1431 297 1863 351
<< fillblock >>
rect 1134 2052 2106 2862
rect 0 1080 3240 2052
rect 1134 216 2106 1080
<< labels >>
flabel locali s 2511 2403 2700 2511 0 FreeSans 240 0 0 0 A
port 1 nsew signal input
flabel locali s 540 567 729 675 0 FreeSans 240 0 0 0 B
port 2 nsew signal input
flabel locali s 2376 2160 2565 2268 0 FreeSans 240 0 0 0 Y
port 3 nsew signal output
flabel metal1 s 2646 405 2835 513 0 FreeSans 240 0 0 0 VPWR
port 4 nsew power bidirectional
flabel metal1 s 189 216 297 378 0 FreeSans 240 0 0 0 VGND
port 5 nsew ground bidirectional
<< end >>
