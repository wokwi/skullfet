magic
tech sky130A
timestamp 1698409033
<< nwell >>
rect 65 50 585 620
<< pwell >>
rect 65 865 585 1380
<< nmos >>
rect 125 1171 530 1211
<< pmos >>
rect 125 245 530 285
<< ndiff >>
rect 233 1320 449 1347
rect 206 1293 449 1320
rect 152 1285 503 1293
rect 152 1255 160 1285
rect 180 1255 503 1285
rect 152 1239 503 1255
rect 125 1211 530 1239
rect 125 1145 530 1171
rect 125 1115 130 1145
rect 150 1131 530 1145
rect 150 1115 206 1131
rect 125 1104 206 1115
rect 125 1077 179 1104
rect 152 1050 179 1077
rect 287 1050 368 1131
rect 449 1104 530 1131
rect 476 1077 530 1104
rect 476 1050 503 1077
rect 152 1023 206 1050
rect 260 1023 395 1050
rect 449 1023 503 1050
rect 152 996 314 1023
rect 341 996 476 1023
rect 206 969 287 996
rect 368 969 476 996
rect 233 915 422 969
rect 233 888 260 915
rect 287 888 314 915
rect 341 888 368 915
rect 395 888 422 915
<< pdiff >>
rect 233 537 260 564
rect 287 537 314 564
rect 341 537 368 564
rect 395 537 422 564
rect 233 483 422 537
rect 206 456 287 483
rect 368 456 476 483
rect 152 429 314 456
rect 341 429 476 456
rect 152 402 206 429
rect 260 402 395 429
rect 449 402 503 429
rect 152 375 179 402
rect 125 348 179 375
rect 125 335 206 348
rect 125 305 130 335
rect 160 321 206 335
rect 287 321 368 402
rect 476 375 503 402
rect 476 348 530 375
rect 449 321 530 348
rect 160 305 530 321
rect 125 285 530 305
rect 125 213 530 245
rect 152 195 503 213
rect 152 165 160 195
rect 180 165 503 195
rect 152 159 503 165
rect 206 132 449 159
rect 233 105 449 132
<< ndiffc >>
rect 160 1255 180 1285
rect 130 1115 150 1145
<< pdiffc >>
rect 130 305 160 335
rect 160 165 180 195
<< psubdiff >>
rect 90 1365 170 1370
rect 90 1325 105 1365
rect 155 1325 170 1365
rect 90 1320 170 1325
<< nsubdiff >>
rect 95 125 165 130
rect 95 90 110 125
rect 150 90 165 125
rect 95 85 165 90
<< psubdiffcont >>
rect 105 1325 155 1365
<< nsubdiffcont >>
rect 110 90 150 125
<< poly >>
rect 10 1171 125 1211
rect 530 1171 660 1211
rect 610 965 660 1171
rect 610 915 620 965
rect 650 915 660 965
rect 610 525 660 915
rect 610 475 620 525
rect 650 475 660 525
rect 610 285 660 475
rect 10 245 125 285
rect 530 245 660 285
<< polycont >>
rect 620 915 650 965
rect 620 475 650 525
<< locali >>
rect 90 1365 170 1370
rect 90 1325 105 1365
rect 155 1325 170 1365
rect 90 1295 170 1325
rect 70 1285 190 1295
rect 70 1260 80 1285
rect 105 1260 160 1285
rect 70 1255 160 1260
rect 180 1255 190 1285
rect 70 1245 190 1255
rect 10 1145 160 1155
rect 10 1115 130 1145
rect 150 1115 160 1145
rect 10 1105 160 1115
rect 10 780 60 1105
rect 10 700 20 780
rect 50 700 60 780
rect 10 345 60 700
rect 610 965 660 985
rect 610 915 620 965
rect 650 915 660 965
rect 610 780 660 915
rect 610 700 620 780
rect 650 700 660 780
rect 610 525 660 700
rect 610 475 620 525
rect 650 475 660 525
rect 610 445 660 475
rect 10 335 170 345
rect 10 305 130 335
rect 160 305 170 335
rect 10 295 170 305
rect 100 195 190 205
rect 100 185 160 195
rect 100 165 105 185
rect 130 165 160 185
rect 180 165 190 195
rect 100 155 190 165
rect 95 125 165 155
rect 95 90 110 125
rect 150 90 165 125
rect 95 85 165 90
<< viali >>
rect 80 1260 105 1285
rect 20 700 50 780
rect 620 700 650 780
rect 105 165 130 185
<< metal1 >>
rect 10 1425 50 1430
rect 10 1385 15 1425
rect 45 1385 50 1425
rect 10 1295 50 1385
rect 233 1320 449 1347
rect 10 1285 110 1295
rect 206 1293 449 1320
rect 10 1260 80 1285
rect 105 1260 110 1285
rect 10 1250 110 1260
rect 152 1239 503 1293
rect 125 1131 530 1239
rect 125 1104 206 1131
rect 125 1077 179 1104
rect 152 1050 179 1077
rect 287 1050 368 1131
rect 449 1104 530 1131
rect 476 1077 530 1104
rect 476 1050 503 1077
rect 152 1023 206 1050
rect 260 1023 395 1050
rect 449 1023 503 1050
rect 152 996 314 1023
rect 341 996 476 1023
rect 206 969 287 996
rect 368 969 476 996
rect 233 915 422 969
rect 71 888 152 915
rect 233 888 260 915
rect 287 888 314 915
rect 341 888 368 915
rect 395 888 422 915
rect 503 888 584 915
rect 44 834 179 888
rect 476 834 611 888
rect 71 807 233 834
rect 422 807 584 834
rect 10 780 62 789
rect 152 780 260 807
rect 395 780 503 807
rect 610 780 660 789
rect 10 700 20 780
rect 50 700 62 780
rect 206 753 314 780
rect 341 753 449 780
rect 10 690 62 700
rect 260 699 395 753
rect 610 700 620 780
rect 650 700 660 780
rect 206 672 314 699
rect 341 672 449 699
rect 610 690 660 700
rect 71 645 260 672
rect 395 645 611 672
rect 44 618 206 645
rect 449 618 611 645
rect 44 591 152 618
rect 503 591 611 618
rect 44 564 125 591
rect 530 564 611 591
rect 71 537 98 564
rect 233 537 260 564
rect 287 537 314 564
rect 341 537 368 564
rect 395 537 422 564
rect 557 537 584 564
rect 233 483 422 537
rect 206 456 287 483
rect 368 456 476 483
rect 152 429 314 456
rect 341 429 476 456
rect 152 402 206 429
rect 260 402 395 429
rect 449 402 503 429
rect 152 375 179 402
rect 125 348 179 375
rect 125 321 206 348
rect 287 321 368 402
rect 476 375 503 402
rect 476 348 530 375
rect 449 321 530 348
rect 125 213 530 321
rect 10 185 135 195
rect 10 165 105 185
rect 130 165 135 185
rect 10 155 135 165
rect 152 159 503 213
rect 10 45 60 155
rect 206 132 449 159
rect 233 105 449 132
rect 10 5 15 45
rect 55 5 60 45
rect 10 0 60 5
<< via1 >>
rect 15 1385 45 1425
rect 15 5 55 45
<< metal2 >>
rect 10 1425 50 1430
rect 10 1385 15 1425
rect 45 1385 50 1425
rect 10 1380 50 1385
rect 233 1320 449 1347
rect 206 1293 449 1320
rect 152 1239 503 1293
rect 125 1131 530 1239
rect 125 1104 206 1131
rect 125 1077 179 1104
rect 152 1050 179 1077
rect 287 1050 368 1131
rect 449 1104 530 1131
rect 476 1077 530 1104
rect 476 1050 503 1077
rect 152 1023 206 1050
rect 260 1023 395 1050
rect 449 1023 503 1050
rect 152 996 314 1023
rect 341 996 476 1023
rect 206 969 287 996
rect 368 969 476 996
rect 233 915 422 969
rect 71 888 152 915
rect 233 888 260 915
rect 287 888 314 915
rect 341 888 368 915
rect 395 888 422 915
rect 503 888 584 915
rect 44 834 179 888
rect 476 834 611 888
rect 71 807 233 834
rect 422 807 584 834
rect 152 780 260 807
rect 395 780 503 807
rect 206 753 314 780
rect 341 753 449 780
rect 260 699 395 753
rect 206 672 314 699
rect 341 672 449 699
rect 71 645 260 672
rect 395 645 611 672
rect 44 618 206 645
rect 449 618 611 645
rect 44 591 152 618
rect 503 591 611 618
rect 44 564 125 591
rect 530 564 611 591
rect 71 537 98 564
rect 233 537 260 564
rect 287 537 314 564
rect 341 537 368 564
rect 395 537 422 564
rect 557 537 584 564
rect 233 483 422 537
rect 206 456 287 483
rect 368 456 476 483
rect 152 429 314 456
rect 341 429 476 456
rect 152 402 206 429
rect 260 402 395 429
rect 449 402 503 429
rect 152 375 179 402
rect 125 348 179 375
rect 125 321 206 348
rect 287 321 368 402
rect 476 375 503 402
rect 476 348 530 375
rect 449 321 530 348
rect 125 213 530 321
rect 152 159 503 213
rect 206 132 449 159
rect 233 105 449 132
rect 10 45 60 50
rect 10 5 15 45
rect 55 5 60 45
rect 10 0 60 5
<< via2 >>
rect 15 1385 45 1425
rect 15 5 55 45
<< metal3 >>
rect 0 1380 670 1430
rect 0 0 670 50 0
<< obsm3 >>
rect 0 90 670 1340
<< fillblock >>
rect 0 0 670 1430
<< labels >>
flabel metal3 s 0 1380 670 1430 0 FreeSans 240 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal3 s 0 0 670 50 0 FreeSans 240 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal1 s 10 695 60 775 0 FreeSans 340 0 0 0 Y
port 3 s signal output
flabel metal1 s 610 695 660 775 0 FreeSans 340 0 0 0 A
port 4 e signal input
<< end >>
