magic
tech sky130A
magscale 1 2
timestamp 1698611668
<< nwell >>
rect 2187 1269 3240 2025
rect 1134 1053 3240 1269
rect 1134 216 2106 1053
<< nmos >>
rect 1215 2403 2025 2511
rect 351 1161 459 1971
<< pmos >>
rect 2781 1161 2889 1971
rect 1215 567 2025 675
<< ndiff >>
rect 1431 2727 1863 2781
rect 1377 2673 1863 2727
rect 1269 2646 1971 2673
rect 1269 2592 1296 2646
rect 1350 2592 1971 2646
rect 1269 2565 1971 2592
rect 1215 2511 2025 2565
rect 1215 2349 2025 2403
rect 1215 2295 1377 2349
rect 1215 2241 1323 2295
rect 1269 2187 1323 2241
rect 1539 2187 1701 2349
rect 1863 2295 1944 2349
rect 1998 2295 2025 2349
rect 1917 2241 2025 2295
rect 1917 2187 1971 2241
rect 1269 2133 1377 2187
rect 1485 2133 1755 2187
rect 1863 2133 1971 2187
rect 1269 2079 1593 2133
rect 1647 2079 1917 2133
rect 1377 2025 1539 2079
rect 1701 2025 1917 2079
rect 297 1917 351 1971
rect 189 1809 351 1917
rect 81 1377 351 1809
rect 135 1323 351 1377
rect 189 1296 351 1323
rect 189 1242 216 1296
rect 270 1242 351 1296
rect 189 1215 351 1242
rect 297 1161 351 1215
rect 459 1944 621 1971
rect 459 1890 513 1944
rect 567 1917 621 1944
rect 1431 1917 1809 2025
rect 567 1890 729 1917
rect 459 1863 729 1890
rect 1431 1863 1485 1917
rect 1539 1863 1593 1917
rect 1647 1863 1701 1917
rect 1755 1863 1809 1917
rect 459 1809 567 1863
rect 675 1809 837 1863
rect 459 1647 513 1809
rect 729 1755 837 1809
rect 729 1701 999 1755
rect 675 1647 945 1701
rect 459 1593 783 1647
rect 837 1593 999 1647
rect 459 1539 729 1593
rect 837 1539 945 1593
rect 459 1485 783 1539
rect 837 1485 999 1539
rect 459 1323 513 1485
rect 675 1431 945 1485
rect 729 1377 999 1431
rect 729 1323 837 1377
rect 459 1269 567 1323
rect 675 1269 783 1323
rect 459 1215 783 1269
rect 459 1161 621 1215
<< pdiff >>
rect 2619 1944 2781 1971
rect 2619 1917 2673 1944
rect 2457 1890 2673 1917
rect 2727 1890 2781 1944
rect 2457 1863 2781 1890
rect 2457 1809 2565 1863
rect 2673 1809 2781 1863
rect 2403 1755 2511 1809
rect 2241 1701 2511 1755
rect 2295 1647 2565 1701
rect 2727 1647 2781 1809
rect 2241 1593 2403 1647
rect 2457 1593 2781 1647
rect 2295 1539 2403 1593
rect 2511 1539 2781 1593
rect 2241 1485 2403 1539
rect 2457 1485 2781 1539
rect 2295 1431 2565 1485
rect 2241 1377 2511 1431
rect 2403 1323 2511 1377
rect 2727 1323 2781 1485
rect 2403 1269 2565 1323
rect 2673 1269 2781 1323
rect 2511 1215 2781 1269
rect 1431 1161 1485 1215
rect 1539 1161 1593 1215
rect 1647 1161 1701 1215
rect 1755 1161 1809 1215
rect 2619 1161 2781 1215
rect 2889 1917 2943 1971
rect 2889 1809 3051 1917
rect 2889 1755 3105 1809
rect 2889 1323 3159 1755
rect 2889 1296 3051 1323
rect 2889 1242 2970 1296
rect 3024 1242 3051 1296
rect 2889 1215 3051 1242
rect 2889 1161 2943 1215
rect 1431 1053 1809 1161
rect 1377 999 1539 1053
rect 1701 999 1917 1053
rect 1269 945 1593 999
rect 1647 945 1917 999
rect 1269 891 1377 945
rect 1485 891 1755 945
rect 1863 891 1971 945
rect 1269 837 1323 891
rect 1215 783 1323 837
rect 1215 729 1377 783
rect 1539 729 1701 891
rect 1917 837 1971 891
rect 1917 783 2025 837
rect 1863 729 1944 783
rect 1998 729 2025 783
rect 1215 675 2025 729
rect 1215 513 2025 567
rect 1269 486 1971 513
rect 1269 432 1890 486
rect 1944 432 1971 486
rect 1269 405 1971 432
rect 1377 351 1863 405
rect 1431 297 1863 351
<< ndiffc >>
rect 1296 2592 1350 2646
rect 1944 2295 1998 2349
rect 216 1242 270 1296
rect 513 1890 567 1944
<< pdiffc >>
rect 2673 1890 2727 1944
rect 2970 1242 3024 1296
rect 1944 729 1998 783
rect 1890 432 1944 486
<< psubdiff >>
rect 27 1242 135 1269
rect 27 1161 81 1242
rect 27 1134 135 1161
<< nsubdiff >>
rect 3105 1242 3186 1269
rect 3159 1161 3186 1242
rect 3105 1107 3186 1161
rect 1917 297 1944 351
rect 2025 297 2052 351
rect 1917 270 2052 297
<< psubdiffcont >>
rect 81 1161 135 1242
<< nsubdiffcont >>
rect 3105 1161 3159 1242
rect 1944 297 2025 351
<< poly >>
rect 1053 2403 1215 2511
rect 2025 2495 2889 2511
rect 2025 2419 2365 2495
rect 2441 2419 2797 2495
rect 2873 2419 2889 2495
rect 2025 2403 2889 2419
rect 351 1971 459 2133
rect 2781 1971 2889 2403
rect 351 675 459 1161
rect 2781 999 2889 1161
rect 351 659 1215 675
rect 351 583 367 659
rect 443 583 799 659
rect 875 583 1215 659
rect 351 567 1215 583
rect 2025 567 2187 675
<< polycont >>
rect 2365 2419 2441 2495
rect 2797 2419 2873 2495
rect 367 583 443 659
rect 799 583 875 659
<< locali >>
rect 1026 2659 1350 2673
rect 1026 2579 1040 2659
rect 1120 2646 1350 2659
rect 1120 2592 1296 2646
rect 1120 2579 1350 2592
rect 1026 2565 1350 2579
rect 2349 2496 2889 2511
rect 2349 2418 2364 2496
rect 2442 2418 2796 2496
rect 2874 2418 2889 2496
rect 2349 2403 2889 2418
rect 1944 2362 2214 2376
rect 1944 2349 2120 2362
rect 1998 2295 2120 2349
rect 1944 2282 2120 2295
rect 2200 2282 2214 2362
rect 1944 2268 2214 2282
rect 486 2146 594 2160
rect 486 2066 500 2146
rect 580 2066 594 2146
rect 486 1944 594 2066
rect 486 1890 513 1944
rect 567 1890 594 1944
rect 2646 2146 2754 2160
rect 2646 2066 2660 2146
rect 2740 2066 2754 2146
rect 2646 1944 2754 2066
rect 2646 1890 2673 1944
rect 2727 1890 2754 1944
rect 81 1242 216 1296
rect 270 1242 297 1296
rect 135 1161 297 1242
rect 81 1026 297 1161
rect 189 1020 297 1026
rect 189 940 200 1020
rect 280 940 297 1020
rect 2943 1242 2970 1296
rect 3024 1269 3051 1296
rect 3024 1242 3159 1269
rect 2943 1161 3105 1242
rect 2943 1053 3159 1161
rect 2943 1039 3051 1053
rect 2943 959 2957 1039
rect 3037 959 3051 1039
rect 2943 945 3051 959
rect 189 920 297 940
rect 1944 796 2214 810
rect 1944 783 2120 796
rect 1998 729 2120 783
rect 1944 716 2120 729
rect 2200 716 2214 796
rect 1944 702 2214 716
rect 351 660 891 675
rect 351 582 366 660
rect 444 582 798 660
rect 876 582 891 660
rect 351 567 891 582
rect 1890 499 2214 513
rect 1890 486 2120 499
rect 1944 432 2120 486
rect 1890 419 2120 432
rect 2200 419 2214 499
rect 1890 405 2214 419
rect 1890 351 2079 405
rect 1890 297 1944 351
rect 2025 297 2079 351
<< viali >>
rect 1040 2579 1120 2659
rect 2364 2495 2442 2496
rect 2364 2419 2365 2495
rect 2365 2419 2441 2495
rect 2441 2419 2442 2495
rect 2364 2418 2442 2419
rect 2796 2495 2874 2496
rect 2796 2419 2797 2495
rect 2797 2419 2873 2495
rect 2873 2419 2874 2495
rect 2796 2418 2874 2419
rect 2120 2282 2200 2362
rect 500 2066 580 2146
rect 2660 2066 2740 2146
rect 200 940 280 1020
rect 2957 959 3037 1039
rect 2120 716 2200 796
rect 366 659 444 660
rect 366 583 367 659
rect 367 583 443 659
rect 443 583 444 659
rect 366 582 444 583
rect 798 659 876 660
rect 798 583 799 659
rect 799 583 875 659
rect 875 583 876 659
rect 798 582 876 583
rect 2120 419 2200 499
<< metal1 >>
rect 1431 2727 1863 2781
rect 1377 2673 1863 2727
rect 486 2659 1134 2673
rect 486 2579 1040 2659
rect 1120 2579 1134 2659
rect 486 2565 1134 2579
rect 1269 2565 1971 2673
rect 486 2146 594 2565
rect 1215 2349 2025 2565
rect 2349 2496 2889 2511
rect 2349 2418 2364 2496
rect 2442 2418 2796 2496
rect 2874 2418 2889 2496
rect 2349 2403 2889 2418
rect 1215 2295 1377 2349
rect 1215 2241 1323 2295
rect 486 2066 500 2146
rect 580 2066 594 2146
rect 1269 2187 1323 2241
rect 1539 2187 1701 2349
rect 1863 2295 2025 2349
rect 1917 2241 2025 2295
rect 2106 2362 2295 2376
rect 2106 2282 2120 2362
rect 2200 2282 2295 2362
rect 2106 2268 2295 2282
rect 1917 2187 1971 2241
rect 1269 2133 1377 2187
rect 1485 2133 1755 2187
rect 1863 2133 1971 2187
rect 2187 2160 2754 2268
rect 2646 2146 2754 2160
rect 1269 2079 1593 2133
rect 1647 2079 1917 2133
rect 486 2052 594 2066
rect 1377 2025 1539 2079
rect 1701 2025 1917 2079
rect 2646 2066 2660 2146
rect 2740 2066 2754 2146
rect 297 1917 621 1971
rect 1431 1917 1809 2025
rect 2646 1971 2754 2066
rect 2619 1917 2943 1971
rect 189 1863 729 1917
rect 1107 1863 1269 1917
rect 1431 1863 1485 1917
rect 1539 1863 1593 1917
rect 1647 1863 1701 1917
rect 1755 1863 1809 1917
rect 1971 1863 2133 1917
rect 2457 1863 3051 1917
rect 189 1809 567 1863
rect 675 1809 837 1863
rect 81 1647 513 1809
rect 729 1755 837 1809
rect 1053 1755 1323 1863
rect 1917 1755 2187 1863
rect 2457 1809 2565 1863
rect 2673 1809 3051 1863
rect 2403 1755 2511 1809
rect 729 1701 999 1755
rect 1107 1701 1431 1755
rect 1809 1701 2133 1755
rect 2241 1701 2511 1755
rect 2727 1755 3105 1809
rect 675 1647 945 1701
rect 1269 1647 1485 1701
rect 1755 1647 1971 1701
rect 2295 1647 2565 1701
rect 2727 1647 3159 1755
rect 81 1593 783 1647
rect 837 1593 999 1647
rect 1377 1593 1593 1647
rect 1647 1593 1863 1647
rect 2241 1593 2403 1647
rect 2457 1593 3159 1647
rect 81 1539 729 1593
rect 837 1539 945 1593
rect 81 1485 783 1539
rect 837 1485 999 1539
rect 1485 1485 1755 1593
rect 2295 1539 2403 1593
rect 2511 1539 3159 1593
rect 2241 1485 2403 1539
rect 2457 1485 3159 1539
rect 81 1377 513 1485
rect 675 1431 945 1485
rect 1377 1431 1593 1485
rect 1647 1431 1863 1485
rect 2295 1431 2565 1485
rect 135 1323 513 1377
rect 729 1377 999 1431
rect 1107 1377 1485 1431
rect 1755 1377 2187 1431
rect 2241 1377 2511 1431
rect 729 1323 837 1377
rect 1053 1323 1377 1377
rect 1863 1323 2187 1377
rect 189 1269 567 1323
rect 675 1269 783 1323
rect 189 1215 783 1269
rect 1053 1269 1269 1323
rect 1971 1269 2187 1323
rect 2403 1323 2511 1377
rect 2727 1323 3159 1485
rect 2403 1269 2565 1323
rect 2673 1269 3051 1323
rect 1053 1215 1215 1269
rect 2025 1215 2187 1269
rect 2511 1215 3051 1269
rect 297 1161 621 1215
rect 1107 1161 1161 1215
rect 1431 1161 1485 1215
rect 1539 1161 1593 1215
rect 1647 1161 1701 1215
rect 1755 1161 1809 1215
rect 2079 1161 2133 1215
rect 2619 1161 2943 1215
rect 1431 1053 1809 1161
rect 180 1030 300 1040
rect 180 930 190 1030
rect 290 930 300 1030
rect 1377 999 1539 1053
rect 1701 999 1917 1053
rect 180 920 300 930
rect 1269 945 1593 999
rect 1647 945 1917 999
rect 1269 891 1377 945
rect 1485 891 1755 945
rect 1863 891 1971 945
rect 1269 837 1323 891
rect 1215 783 1323 837
rect 1215 729 1377 783
rect 1539 729 1701 891
rect 1917 837 1971 891
rect 1917 783 2025 837
rect 2646 810 2754 1161
rect 1863 729 2025 783
rect 351 660 891 675
rect 351 582 366 660
rect 444 582 798 660
rect 876 582 891 660
rect 351 567 891 582
rect 1215 513 2025 729
rect 2106 796 2754 810
rect 2106 716 2120 796
rect 2200 716 2754 796
rect 2106 702 2754 716
rect 2943 1039 3051 1053
rect 2943 959 2957 1039
rect 3037 959 3051 1039
rect 2943 513 3051 959
rect 1269 405 1971 513
rect 2106 503 3051 513
rect 2106 499 2953 503
rect 2106 419 2120 499
rect 2200 419 2953 499
rect 2106 415 2953 419
rect 3041 415 3051 503
rect 2106 405 3051 415
rect 1377 351 1863 405
rect 1431 297 1863 351
<< via1 >>
rect 190 1020 290 1030
rect 190 940 200 1020
rect 200 940 280 1020
rect 280 940 290 1020
rect 190 930 290 940
rect 2953 415 3041 503
<< metal2 >>
rect 1431 2727 1863 2781
rect 1377 2673 1863 2727
rect 1269 2565 1971 2673
rect 1215 2349 2025 2565
rect 1215 2295 1377 2349
rect 1215 2241 1323 2295
rect 1269 2187 1323 2241
rect 1539 2187 1701 2349
rect 1863 2295 2025 2349
rect 1917 2241 2025 2295
rect 1917 2187 1971 2241
rect 1269 2133 1377 2187
rect 1485 2133 1755 2187
rect 1863 2133 1971 2187
rect 1269 2079 1593 2133
rect 1647 2079 1917 2133
rect 1377 2025 1539 2079
rect 1701 2025 1917 2079
rect 297 1917 621 1971
rect 1431 1917 1809 2025
rect 2619 1917 2943 1971
rect 189 1863 729 1917
rect 1431 1863 1485 1917
rect 1539 1863 1593 1917
rect 1647 1863 1701 1917
rect 1755 1863 1809 1917
rect 2457 1863 3051 1917
rect 189 1809 567 1863
rect 675 1809 837 1863
rect 2457 1809 2565 1863
rect 2673 1809 3051 1863
rect 81 1647 513 1809
rect 729 1755 837 1809
rect 2403 1755 2511 1809
rect 729 1701 999 1755
rect 2241 1701 2511 1755
rect 2727 1755 3105 1809
rect 675 1647 945 1701
rect 2295 1647 2565 1701
rect 2727 1647 3159 1755
rect 81 1593 783 1647
rect 837 1593 999 1647
rect 2241 1593 2403 1647
rect 2457 1593 3159 1647
rect 81 1539 729 1593
rect 837 1539 945 1593
rect 2295 1539 2403 1593
rect 2511 1539 3159 1593
rect 81 1485 783 1539
rect 837 1485 999 1539
rect 2241 1485 2403 1539
rect 2457 1485 3159 1539
rect 81 1377 513 1485
rect 675 1431 945 1485
rect 2295 1431 2565 1485
rect 135 1323 513 1377
rect 729 1377 999 1431
rect 2241 1377 2511 1431
rect 729 1323 837 1377
rect 2403 1323 2511 1377
rect 2727 1323 3159 1485
rect 189 1269 567 1323
rect 675 1269 783 1323
rect 2403 1269 2565 1323
rect 2673 1269 3051 1323
rect 189 1215 783 1269
rect 2511 1215 3051 1269
rect 297 1161 621 1215
rect 1431 1161 1485 1215
rect 1539 1161 1593 1215
rect 1647 1161 1701 1215
rect 1755 1161 1809 1215
rect 2619 1161 2943 1215
rect 1431 1053 1809 1161
rect 180 1030 300 1040
rect 180 930 190 1030
rect 290 930 300 1030
rect 1377 999 1539 1053
rect 1701 999 1917 1053
rect 180 210 300 930
rect 1269 945 1593 999
rect 1647 945 1917 999
rect 1269 891 1377 945
rect 1485 891 1755 945
rect 1863 891 1971 945
rect 1269 837 1323 891
rect 1215 783 1323 837
rect 1215 729 1377 783
rect 1539 729 1701 891
rect 1917 837 1971 891
rect 1917 783 2025 837
rect 1863 729 2025 783
rect 1215 513 2025 729
rect 1269 405 1971 513
rect 2940 503 3060 520
rect 2940 415 2953 503
rect 3041 415 3060 503
rect 1377 351 1863 405
rect 1431 297 1863 351
rect 180 150 190 210
rect 290 150 300 210
rect 180 140 300 150
rect 2940 70 3060 415
rect 2940 10 2950 70
rect 3050 10 3060 70
rect 2940 0 3060 10
<< via2 >>
rect 190 150 290 210
rect 2950 10 3050 70
<< metal3 >>
rect 0 210 3240 220
rect 0 150 190 210
rect 290 150 3240 210
rect 0 140 3240 150
rect 0 70 3240 80
rect 0 10 2950 70
rect 3050 10 3240 70
rect 0 0 3240 10
<< fillblock >>
rect 1134 2052 2106 2862
rect 0 1080 3240 2052
rect 1134 216 2106 1080
<< labels >>
flabel metal1 s 2349 2403 2889 2511 0 FreeSans 240 0 0 0 A
port 1 nsew signal input
flabel metal1 s 351 567 891 675 0 FreeSans 240 0 0 0 B
port 2 nsew signal input
flabel metal1 s 2187 2160 2754 2268 0 FreeSans 240 0 0 0 Y
port 3 nsew signal output
flabel metal3 s 0 0 3240 80 0 FreeSans 240 0 0 0 VPWR
port 4 nsew power input
flabel metal3 s 0 140 3240 220 0 FreeSans 240 0 0 0 VGND
port 5 nsew ground input
<< end >>
