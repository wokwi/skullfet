magic
tech sky130A
timestamp 1641001583
<< nwell >>
rect 3050 600 8250 6300
<< pwell >>
rect 3050 8750 8250 13900
<< nmos >>
rect 3650 11810 7700 12210
<< pmos >>
rect 3650 2550 7700 2950
<< ndiff >>
rect 4730 13300 6890 13570
rect 4460 13030 6890 13300
rect 3920 12950 7430 13030
rect 3920 12650 4000 12950
rect 4200 12650 7430 12950
rect 3920 12490 7430 12650
rect 3650 12210 7700 12490
rect 3650 11550 7700 11810
rect 3650 11250 3700 11550
rect 3900 11410 7700 11550
rect 3900 11250 4460 11410
rect 3650 11140 4460 11250
rect 3650 10870 4190 11140
rect 3920 10600 4190 10870
rect 5270 10600 6080 11410
rect 6890 11140 7700 11410
rect 7160 10870 7700 11140
rect 7160 10600 7430 10870
rect 3920 10330 4460 10600
rect 5000 10330 6350 10600
rect 6890 10330 7430 10600
rect 3920 10060 5540 10330
rect 5810 10060 7160 10330
rect 4460 9790 5270 10060
rect 6080 9790 7160 10060
rect 4730 9250 6620 9790
rect 4730 8980 5000 9250
rect 5270 8980 5540 9250
rect 5810 8980 6080 9250
rect 6350 8980 6620 9250
<< pdiff >>
rect 4730 5470 5000 5740
rect 5270 5470 5540 5740
rect 5810 5470 6080 5740
rect 6350 5470 6620 5740
rect 4730 4930 6620 5470
rect 4460 4660 5270 4930
rect 6080 4660 7160 4930
rect 3920 4390 5540 4660
rect 5810 4390 7160 4660
rect 3920 4120 4460 4390
rect 5000 4120 6350 4390
rect 6890 4120 7430 4390
rect 3920 3850 4190 4120
rect 3650 3580 4190 3850
rect 3650 3450 4460 3580
rect 3650 3150 3700 3450
rect 4000 3310 4460 3450
rect 5270 3310 6080 4120
rect 7160 3850 7430 4120
rect 7160 3580 7700 3850
rect 6890 3310 7700 3580
rect 4000 3150 7700 3310
rect 3650 2950 7700 3150
rect 3650 2230 7700 2550
rect 3920 2050 7430 2230
rect 3920 1750 4000 2050
rect 4200 1750 7430 2050
rect 3920 1690 7430 1750
rect 4460 1420 6890 1690
rect 4730 1150 6890 1420
<< ndiffc >>
rect 4000 12650 4200 12950
rect 3700 11250 3900 11550
<< pdiffc >>
rect 3700 3150 4000 3450
rect 4000 1750 4200 2050
<< psubdiff >>
rect 3300 13750 4400 13800
rect 3300 13350 3450 13750
rect 3950 13700 4400 13750
rect 3950 13500 4000 13700
rect 4300 13500 4400 13700
rect 7100 13700 7500 13800
rect 3950 13400 4400 13500
rect 3950 13350 4100 13400
rect 3300 13300 4100 13350
rect 7100 13500 7200 13700
rect 7400 13500 7500 13700
rect 7100 13400 7500 13500
rect 4700 11100 5100 11200
rect 4700 10900 4800 11100
rect 5000 10900 5100 11100
rect 4700 10800 5100 10900
rect 6300 11100 6700 11200
rect 6300 10900 6400 11100
rect 6600 10900 6700 11100
rect 6300 10800 6700 10900
rect 5500 8850 5850 8900
rect 5500 8800 5550 8850
rect 5800 8800 5850 8850
rect 5500 8750 5850 8800
<< nsubdiff >>
rect 5500 6100 5900 6200
rect 5500 6000 5600 6100
rect 5800 6000 5900 6100
rect 5500 5900 5900 6000
rect 4600 3800 5000 3900
rect 4600 3600 4700 3800
rect 4900 3600 5000 3800
rect 4600 3500 5000 3600
rect 6300 3800 6700 3900
rect 6300 3600 6400 3800
rect 6600 3600 6700 3800
rect 6300 3500 6700 3600
rect 3350 1350 4050 1400
rect 3350 1100 3500 1350
rect 3900 1300 4050 1350
rect 3900 1200 4400 1300
rect 3900 1100 4000 1200
rect 4300 1100 4400 1200
rect 7100 1400 7700 1500
rect 3350 1000 4400 1100
rect 7100 1000 7200 1400
rect 7600 1000 7700 1400
rect 7100 900 7700 1000
<< psubdiffcont >>
rect 3450 13350 3950 13750
rect 4000 13500 4300 13700
rect 7200 13500 7400 13700
rect 4800 10900 5000 11100
rect 6400 10900 6600 11100
rect 5550 8800 5800 8850
<< nsubdiffcont >>
rect 5600 6000 5800 6100
rect 4700 3600 4900 3800
rect 6400 3600 6600 3800
rect 3500 1100 3900 1350
rect 4000 1100 4300 1200
rect 7200 1000 7600 1400
<< poly >>
rect 2500 11810 3650 12210
rect 7700 11810 9000 12210
rect 8500 9750 9000 11810
rect 8500 9250 8600 9750
rect 8900 9250 9000 9750
rect 8500 5350 9000 9250
rect 8500 4850 8600 5350
rect 8900 4850 9000 5350
rect 8500 2950 9000 4850
rect 2500 2550 3650 2950
rect 7700 2550 9000 2950
<< polycont >>
rect 8600 9250 8900 9750
rect 8600 4850 8900 5350
<< locali >>
rect 3300 13750 4400 13800
rect 3300 13350 3450 13750
rect 3950 13700 4400 13750
rect 3950 13500 4000 13700
rect 4300 13500 4400 13700
rect 3950 13400 4400 13500
rect 7100 13700 8200 13800
rect 7100 13500 7200 13700
rect 7400 13500 7900 13700
rect 8100 13600 8200 13700
rect 8100 13500 8300 13600
rect 7100 13400 8300 13500
rect 3950 13350 4100 13400
rect 3300 13050 4100 13350
rect 3100 12950 4300 13050
rect 3100 12700 3200 12950
rect 3450 12700 4000 12950
rect 3100 12650 4000 12700
rect 4200 12650 4300 12950
rect 3100 12550 4300 12650
rect 2500 11550 4000 11650
rect 2500 11250 3700 11550
rect 3900 11250 4000 11550
rect 2500 11150 4000 11250
rect 2500 3550 3000 11150
rect 4700 11100 5100 11200
rect 6300 11100 6700 11200
rect 8000 11100 8300 13400
rect 4700 10900 4800 11100
rect 5000 10900 6400 11100
rect 6600 10900 8300 11100
rect 4700 10800 5100 10900
rect 6300 10800 6700 10900
rect 8000 9700 8300 10900
rect 6800 9500 8300 9700
rect 8500 9750 9000 9950
rect 6800 8900 7000 9500
rect 5500 8850 7000 8900
rect 5500 8800 5550 8850
rect 5800 8800 7000 8850
rect 5500 8750 7000 8800
rect 8500 9250 8600 9750
rect 8900 9250 9000 9750
rect 5500 6100 5900 6200
rect 5500 6000 5600 6100
rect 5800 6000 7300 6100
rect 5500 5900 7300 6000
rect 7100 5300 7300 5900
rect 8500 5350 9000 9250
rect 7100 5100 8200 5300
rect 4600 3800 5000 3900
rect 6300 3800 6700 3900
rect 7900 3800 8200 5100
rect 8500 4850 8600 5350
rect 8900 4850 9000 5350
rect 8500 4550 9000 4850
rect 4600 3600 4700 3800
rect 4900 3600 6400 3800
rect 6600 3600 8200 3800
rect 2500 3450 4100 3550
rect 4600 3500 5000 3600
rect 6300 3500 6700 3600
rect 2500 3150 3700 3450
rect 4000 3150 4100 3450
rect 2500 3050 4100 3150
rect 3400 2050 4300 2150
rect 3400 1950 4000 2050
rect 3400 1750 3450 1950
rect 3700 1750 4000 1950
rect 4200 1750 4300 2050
rect 3400 1650 4300 1750
rect 3350 1350 4050 1650
rect 7900 1500 8200 3600
rect 3350 1100 3500 1350
rect 3900 1300 4050 1350
rect 7100 1400 8200 1500
rect 3900 1200 4400 1300
rect 3900 1100 4000 1200
rect 4300 1100 4400 1200
rect 3350 1000 4400 1100
rect 7100 1000 7200 1400
rect 7600 1000 7900 1400
rect 8100 1000 8200 1400
rect 7100 900 8200 1000
<< viali >>
rect 7900 13500 8100 13700
rect 3200 12700 3450 12950
rect 3450 1750 3700 1950
rect 7900 1000 8100 1400
<< metal1 >>
rect 0 14000 10700 14400
rect 2500 13050 2900 14000
rect 7800 13700 8300 14000
rect 4730 13300 6890 13570
rect 7800 13500 7900 13700
rect 8100 13500 8300 13700
rect 7800 13400 8300 13500
rect 2500 12950 3500 13050
rect 4460 13030 6890 13300
rect 2500 12700 3200 12950
rect 3450 12700 3500 12950
rect 2500 12600 3500 12700
rect 3920 12490 7430 13030
rect 3650 11410 7700 12490
rect 3650 11140 4460 11410
rect 3650 10870 4190 11140
rect 3920 10600 4190 10870
rect 5270 10600 6080 11410
rect 6890 11140 7700 11410
rect 7160 10870 7700 11140
rect 7160 10600 7430 10870
rect 3920 10330 4460 10600
rect 5000 10330 6350 10600
rect 6890 10330 7430 10600
rect 3920 10060 5540 10330
rect 5810 10060 7160 10330
rect 4460 9790 5270 10060
rect 6080 9790 7160 10060
rect 4730 9250 6620 9790
rect 3110 8980 3920 9250
rect 4730 8980 5000 9250
rect 5270 8980 5540 9250
rect 5810 8980 6080 9250
rect 6350 8980 6620 9250
rect 7430 8980 8240 9250
rect 2840 8440 4190 8980
rect 7160 8440 8510 8980
rect 3110 8170 4730 8440
rect 6620 8170 8240 8440
rect 3920 7900 5000 8170
rect 6350 7900 7430 8170
rect 4460 7630 5540 7900
rect 5810 7630 6890 7900
rect 5000 7090 6350 7630
rect 4460 6820 5540 7090
rect 5810 6820 6890 7090
rect 3110 6550 5000 6820
rect 6350 6550 8510 6820
rect 2840 6280 4460 6550
rect 6890 6280 8510 6550
rect 2840 6010 3920 6280
rect 7430 6010 8510 6280
rect 2840 5740 3650 6010
rect 7700 5740 8510 6010
rect 3110 5470 3380 5740
rect 4730 5470 5000 5740
rect 5270 5470 5540 5740
rect 5810 5470 6080 5740
rect 6350 5470 6620 5740
rect 7970 5470 8240 5740
rect 4730 4930 6620 5470
rect 4460 4660 5270 4930
rect 6080 4660 7160 4930
rect 3920 4390 5540 4660
rect 5810 4390 7160 4660
rect 3920 4120 4460 4390
rect 5000 4120 6350 4390
rect 6890 4120 7430 4390
rect 3920 3850 4190 4120
rect 3650 3580 4190 3850
rect 3650 3310 4460 3580
rect 5270 3310 6080 4120
rect 7160 3850 7430 4120
rect 7160 3580 7700 3850
rect 6890 3310 7700 3580
rect 3650 2230 7700 3310
rect 2500 1950 3750 2050
rect 2500 1750 3450 1950
rect 3700 1750 3750 1950
rect 2500 1650 3750 1750
rect 3920 1690 7430 2230
rect 2500 400 3000 1650
rect 4460 1420 6890 1690
rect 4730 1150 6890 1420
rect 7700 1400 8200 1500
rect 7700 1000 7900 1400
rect 8100 1000 8200 1400
rect 7700 400 8200 1000
rect 0 0 10700 400
<< metal2 >>
rect 4730 13300 6890 13570
rect 4460 13030 6890 13300
rect 3920 12490 7430 13030
rect 3650 11410 7700 12490
rect 3650 11140 4460 11410
rect 3650 10870 4190 11140
rect 3920 10600 4190 10870
rect 5270 10600 6080 11410
rect 6890 11140 7700 11410
rect 7160 10870 7700 11140
rect 7160 10600 7430 10870
rect 3920 10330 4460 10600
rect 5000 10330 6350 10600
rect 6890 10330 7430 10600
rect 3920 10060 5540 10330
rect 5810 10060 7160 10330
rect 4460 9790 5270 10060
rect 6080 9790 7160 10060
rect 4730 9250 6620 9790
rect 3110 8980 3920 9250
rect 4730 8980 5000 9250
rect 5270 8980 5540 9250
rect 5810 8980 6080 9250
rect 6350 8980 6620 9250
rect 7430 8980 8240 9250
rect 2840 8440 4190 8980
rect 7160 8440 8510 8980
rect 3110 8170 4730 8440
rect 6620 8170 8240 8440
rect 3920 7900 5000 8170
rect 6350 7900 7430 8170
rect 4460 7630 5540 7900
rect 5810 7630 6890 7900
rect 5000 7090 6350 7630
rect 4460 6820 5540 7090
rect 5810 6820 6890 7090
rect 3110 6550 5000 6820
rect 6350 6550 8510 6820
rect 2840 6280 4460 6550
rect 6890 6280 8510 6550
rect 2840 6010 3920 6280
rect 7430 6010 8510 6280
rect 2840 5740 3650 6010
rect 7700 5740 8510 6010
rect 3110 5470 3380 5740
rect 4730 5470 5000 5740
rect 5270 5470 5540 5740
rect 5810 5470 6080 5740
rect 6350 5470 6620 5740
rect 7970 5470 8240 5740
rect 4730 4930 6620 5470
rect 4460 4660 5270 4930
rect 6080 4660 7160 4930
rect 3920 4390 5540 4660
rect 5810 4390 7160 4660
rect 3920 4120 4460 4390
rect 5000 4120 6350 4390
rect 6890 4120 7430 4390
rect 3920 3850 4190 4120
rect 3650 3580 4190 3850
rect 3650 3310 4460 3580
rect 5270 3310 6080 4120
rect 7160 3850 7430 4120
rect 7160 3580 7700 3850
rect 6890 3310 7700 3580
rect 3650 2230 7700 3310
rect 3920 1690 7430 2230
rect 4460 1420 6890 1690
rect 4730 1150 6890 1420
<< metal3 >>
rect 4730 13300 6890 13570
rect 4460 13030 6890 13300
rect 3920 12490 7430 13030
rect 3650 11410 7700 12490
rect 3650 11140 4460 11410
rect 3650 10870 4190 11140
rect 3920 10600 4190 10870
rect 5270 10600 6080 11410
rect 6890 11140 7700 11410
rect 7160 10870 7700 11140
rect 7160 10600 7430 10870
rect 3920 10330 4460 10600
rect 5000 10330 6350 10600
rect 6890 10330 7430 10600
rect 3920 10060 5540 10330
rect 5810 10060 7160 10330
rect 4460 9790 5270 10060
rect 6080 9790 7160 10060
rect 4730 9250 6620 9790
rect 3110 8980 3920 9250
rect 4730 8980 5000 9250
rect 5270 8980 5540 9250
rect 5810 8980 6080 9250
rect 6350 8980 6620 9250
rect 7430 8980 8240 9250
rect 2840 8440 4190 8980
rect 7160 8440 8510 8980
rect 3110 8170 4730 8440
rect 6620 8170 8240 8440
rect 3920 7900 5000 8170
rect 6350 7900 7430 8170
rect 4460 7630 5540 7900
rect 5810 7630 6890 7900
rect 5000 7090 6350 7630
rect 4460 6820 5540 7090
rect 5810 6820 6890 7090
rect 3110 6550 5000 6820
rect 6350 6550 8510 6820
rect 2840 6280 4460 6550
rect 6890 6280 8510 6550
rect 2840 6010 3920 6280
rect 7430 6010 8510 6280
rect 2840 5740 3650 6010
rect 7700 5740 8510 6010
rect 3110 5470 3380 5740
rect 4730 5470 5000 5740
rect 5270 5470 5540 5740
rect 5810 5470 6080 5740
rect 6350 5470 6620 5740
rect 7970 5470 8240 5740
rect 4730 4930 6620 5470
rect 4460 4660 5270 4930
rect 6080 4660 7160 4930
rect 3920 4390 5540 4660
rect 5810 4390 7160 4660
rect 3920 4120 4460 4390
rect 5000 4120 6350 4390
rect 6890 4120 7430 4390
rect 3920 3850 4190 4120
rect 3650 3580 4190 3850
rect 3650 3310 4460 3580
rect 5270 3310 6080 4120
rect 7160 3850 7430 4120
rect 7160 3580 7700 3850
rect 6890 3310 7700 3580
rect 3650 2230 7700 3310
rect 3920 1690 7430 2230
rect 4460 1420 6890 1690
rect 4730 1150 6890 1420
<< metal4 >>
rect 4730 13300 6890 13570
rect 4460 13030 6890 13300
rect 3920 12490 7430 13030
rect 3650 11410 7700 12490
rect 3650 11140 4460 11410
rect 3650 10870 4190 11140
rect 3920 10600 4190 10870
rect 5270 10600 6080 11410
rect 6890 11140 7700 11410
rect 7160 10870 7700 11140
rect 7160 10600 7430 10870
rect 3920 10330 4460 10600
rect 5000 10330 6350 10600
rect 6890 10330 7430 10600
rect 3920 10060 5540 10330
rect 5810 10060 7160 10330
rect 4460 9790 5270 10060
rect 6080 9790 7160 10060
rect 4730 9250 6620 9790
rect 3110 8980 3920 9250
rect 4730 8980 5000 9250
rect 5270 8980 5540 9250
rect 5810 8980 6080 9250
rect 6350 8980 6620 9250
rect 7430 8980 8240 9250
rect 2840 8440 4190 8980
rect 7160 8440 8510 8980
rect 3110 8170 4730 8440
rect 6620 8170 8240 8440
rect 3920 7900 5000 8170
rect 6350 7900 7430 8170
rect 4460 7630 5540 7900
rect 5810 7630 6890 7900
rect 5000 7090 6350 7630
rect 4460 6820 5540 7090
rect 5810 6820 6890 7090
rect 3110 6550 5000 6820
rect 6350 6550 8510 6820
rect 2840 6280 4460 6550
rect 6890 6280 8510 6550
rect 2840 6010 3920 6280
rect 7430 6010 8510 6280
rect 2840 5740 3650 6010
rect 7700 5740 8510 6010
rect 3110 5470 3380 5740
rect 4730 5470 5000 5740
rect 5270 5470 5540 5740
rect 5810 5470 6080 5740
rect 6350 5470 6620 5740
rect 7970 5470 8240 5740
rect 4730 4930 6620 5470
rect 4460 4660 5270 4930
rect 6080 4660 7160 4930
rect 3920 4390 5540 4660
rect 5810 4390 7160 4660
rect 3920 4120 4460 4390
rect 5000 4120 6350 4390
rect 6890 4120 7430 4390
rect 3920 3850 4190 4120
rect 3650 3580 4190 3850
rect 3650 3310 4460 3580
rect 5270 3310 6080 4120
rect 7160 3850 7430 4120
rect 7160 3580 7700 3850
rect 6890 3310 7700 3580
rect 3650 2230 7700 3310
rect 3920 1690 7430 2230
rect 4460 1420 6890 1690
rect 4730 1150 6890 1420
<< metal5 >>
rect 4730 13300 6890 13570
rect 4460 13030 6890 13300
rect 3920 12490 7430 13030
rect 3650 11410 7700 12490
rect 3650 11140 4460 11410
rect 3650 10870 4190 11140
rect 3920 10600 4190 10870
rect 5270 10600 6080 11410
rect 6890 11140 7700 11410
rect 7160 10870 7700 11140
rect 7160 10600 7430 10870
rect 3920 10330 4460 10600
rect 5000 10330 6350 10600
rect 6890 10330 7430 10600
rect 3920 10060 5540 10330
rect 5810 10060 7160 10330
rect 4460 9790 5270 10060
rect 6080 9790 7160 10060
rect 4730 9250 6620 9790
rect 3110 8980 3920 9250
rect 4730 8980 5000 9250
rect 5270 8980 5540 9250
rect 5810 8980 6080 9250
rect 6350 8980 6620 9250
rect 7430 8980 8240 9250
rect 2840 8440 4190 8980
rect 7160 8440 8510 8980
rect 3110 8170 4730 8440
rect 6620 8170 8240 8440
rect 3920 7900 5000 8170
rect 6350 7900 7430 8170
rect 4460 7630 5540 7900
rect 5810 7630 6890 7900
rect 5000 7090 6350 7630
rect 4460 6820 5540 7090
rect 5810 6820 6890 7090
rect 3110 6550 5000 6820
rect 6350 6550 8510 6820
rect 2840 6280 4460 6550
rect 6890 6280 8510 6550
rect 2840 6010 3920 6280
rect 7430 6010 8510 6280
rect 2840 5740 3650 6010
rect 7700 5740 8510 6010
rect 3110 5470 3380 5740
rect 4730 5470 5000 5740
rect 5270 5470 5540 5740
rect 5810 5470 6080 5740
rect 6350 5470 6620 5740
rect 7970 5470 8240 5740
rect 4730 4930 6620 5470
rect 4460 4660 5270 4930
rect 6080 4660 7160 4930
rect 3920 4390 5540 4660
rect 5810 4390 7160 4660
rect 3920 4120 4460 4390
rect 5000 4120 6350 4390
rect 6890 4120 7430 4390
rect 3920 3850 4190 4120
rect 3650 3580 4190 3850
rect 3650 3310 4460 3580
rect 5270 3310 6080 4120
rect 7160 3850 7430 4120
rect 7160 3580 7700 3850
rect 6890 3310 7700 3580
rect 3650 2230 7700 3310
rect 3920 1690 7430 2230
rect 4460 1420 6890 1690
rect 4730 1150 6890 1420
<< labels >>
flabel metal1 s 2500 12600 2900 13050 0 FreeSans 240 90 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 2500 1650 3000 2050 0 FreeSans 240 90 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 2500 7050 3000 7850 0 FreeSans 340 0 0 0 Y
port 3 s signal output
flabel locali s 8500 7050 9000 7850 0 FreeSans 340 0 0 0 A
port 4 e signal input
<< end >>
