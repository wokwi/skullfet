magic
tech sky130A
timestamp 1640345212
<< nwell >>
rect 55 0 575 570
<< pwell >>
rect 55 815 575 1330
<< nmos >>
rect 115 1121 520 1161
<< pmos >>
rect 115 195 520 235
<< ndiff >>
rect 223 1270 439 1297
rect 196 1243 439 1270
rect 142 1235 493 1243
rect 142 1205 150 1235
rect 170 1205 493 1235
rect 142 1189 493 1205
rect 115 1161 520 1189
rect 115 1095 520 1121
rect 115 1065 120 1095
rect 140 1081 520 1095
rect 140 1065 196 1081
rect 115 1054 196 1065
rect 115 1027 169 1054
rect 142 1000 169 1027
rect 277 1000 358 1081
rect 439 1054 520 1081
rect 466 1027 520 1054
rect 466 1000 493 1027
rect 142 973 196 1000
rect 250 973 385 1000
rect 439 973 493 1000
rect 142 946 304 973
rect 331 946 466 973
rect 196 919 277 946
rect 358 919 466 946
rect 223 865 412 919
rect 223 838 250 865
rect 277 838 304 865
rect 331 838 358 865
rect 385 838 412 865
<< pdiff >>
rect 223 487 250 514
rect 277 487 304 514
rect 331 487 358 514
rect 385 487 412 514
rect 223 433 412 487
rect 196 406 277 433
rect 358 406 466 433
rect 142 379 304 406
rect 331 379 466 406
rect 142 352 196 379
rect 250 352 385 379
rect 439 352 493 379
rect 142 325 169 352
rect 115 298 169 325
rect 115 285 196 298
rect 115 255 120 285
rect 150 271 196 285
rect 277 271 358 352
rect 466 325 493 352
rect 466 298 520 325
rect 439 271 520 298
rect 150 255 520 271
rect 115 235 520 255
rect 115 163 520 195
rect 142 145 493 163
rect 142 115 150 145
rect 170 115 493 145
rect 142 109 493 115
rect 196 82 439 109
rect 223 55 439 82
<< ndiffc >>
rect 150 1205 170 1235
rect 120 1065 140 1095
<< pdiffc >>
rect 120 255 150 285
rect 150 115 170 145
<< psubdiff >>
rect 80 1315 160 1320
rect 80 1275 95 1315
rect 145 1275 160 1315
rect 80 1270 160 1275
<< nsubdiff >>
rect 85 75 155 80
rect 85 40 100 75
rect 140 40 155 75
rect 85 35 155 40
<< psubdiffcont >>
rect 95 1275 145 1315
<< nsubdiffcont >>
rect 100 40 140 75
<< poly >>
rect 0 1121 115 1161
rect 520 1121 650 1161
rect 600 915 650 1121
rect 600 865 610 915
rect 640 865 650 915
rect 600 475 650 865
rect 600 425 610 475
rect 640 425 650 475
rect 600 235 650 425
rect 0 195 115 235
rect 520 195 650 235
<< polycont >>
rect 610 865 640 915
rect 610 425 640 475
<< locali >>
rect 80 1315 160 1320
rect 80 1275 95 1315
rect 145 1275 160 1315
rect 80 1245 160 1275
rect 60 1235 180 1245
rect 60 1205 70 1235
rect 100 1205 150 1235
rect 170 1205 180 1235
rect 60 1195 180 1205
rect 0 1095 150 1105
rect 0 1065 120 1095
rect 140 1065 150 1095
rect 0 1055 150 1065
rect 0 295 50 1055
rect 600 915 650 935
rect 600 865 610 915
rect 640 865 650 915
rect 600 475 650 865
rect 600 425 610 475
rect 640 425 650 475
rect 600 395 650 425
rect 0 285 160 295
rect 0 255 120 285
rect 150 255 160 285
rect 0 245 160 255
rect 90 145 180 155
rect 90 115 100 145
rect 130 115 150 145
rect 170 115 180 145
rect 90 105 180 115
rect 85 75 155 105
rect 85 40 100 75
rect 140 40 155 75
rect 85 35 155 40
<< viali >>
rect 70 1205 100 1235
rect 100 115 130 145
<< metal1 >>
rect 0 1235 110 1245
rect 0 1205 70 1235
rect 100 1205 110 1235
rect 0 1195 110 1205
rect 61 838 142 865
rect 493 838 574 865
rect 34 784 169 838
rect 466 784 601 838
rect 61 757 223 784
rect 412 757 574 784
rect 142 730 250 757
rect 385 730 493 757
rect 196 703 304 730
rect 331 703 439 730
rect 250 649 385 703
rect 196 622 304 649
rect 331 622 439 649
rect 61 595 250 622
rect 385 595 601 622
rect 34 568 196 595
rect 439 568 601 595
rect 34 541 142 568
rect 493 541 601 568
rect 34 514 115 541
rect 520 514 601 541
rect 61 487 88 514
rect 547 487 574 514
rect 0 145 140 155
rect 0 115 100 145
rect 130 115 140 145
rect 0 105 140 115
<< labels >>
flabel metal1 s 0 1195 50 1245 0 FreeSans 240 90 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 0 105 50 155 0 FreeSans 240 90 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 0 645 50 725 0 FreeSans 340 0 0 0 Y
port 3 s signal output
flabel locali s 600 645 650 725 0 FreeSans 340 0 0 0 A
port 4 e signal input
flabel metal1 s 60 105 110 155 0 FreeSans 240 90 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 60 1195 110 1245 0 FreeSans 240 90 0 0 VNB
port 6 nsew ground bidirectional
<< end >>
