magic
tech gf180mcuC
timestamp 1669746995
<< nwell >>
rect 305 60 825 630
<< pwell >>
rect 305 875 825 1390
<< nmos >>
rect 365 1181 770 1221
<< pmos >>
rect 365 255 770 295
<< ndiff >>
rect 473 1330 689 1357
rect 446 1303 689 1330
rect 392 1295 743 1303
rect 392 1265 400 1295
rect 420 1265 743 1295
rect 392 1249 743 1265
rect 365 1221 770 1249
rect 365 1155 770 1181
rect 365 1125 370 1155
rect 390 1141 770 1155
rect 390 1125 446 1141
rect 365 1114 446 1125
rect 365 1087 419 1114
rect 392 1060 419 1087
rect 527 1060 608 1141
rect 689 1114 770 1141
rect 716 1087 770 1114
rect 716 1060 743 1087
rect 392 1033 446 1060
rect 500 1033 635 1060
rect 689 1033 743 1060
rect 392 1006 554 1033
rect 581 1006 716 1033
rect 446 979 527 1006
rect 608 979 716 1006
rect 473 925 662 979
rect 473 898 500 925
rect 527 898 554 925
rect 581 898 608 925
rect 635 898 662 925
<< pdiff >>
rect 473 547 500 574
rect 527 547 554 574
rect 581 547 608 574
rect 635 547 662 574
rect 473 493 662 547
rect 446 466 527 493
rect 608 466 716 493
rect 392 439 554 466
rect 581 439 716 466
rect 392 412 446 439
rect 500 412 635 439
rect 689 412 743 439
rect 392 385 419 412
rect 365 358 419 385
rect 365 345 446 358
rect 365 315 370 345
rect 400 331 446 345
rect 527 331 608 412
rect 716 385 743 412
rect 716 358 770 385
rect 689 331 770 358
rect 400 315 770 331
rect 365 295 770 315
rect 365 223 770 255
rect 392 205 743 223
rect 392 175 400 205
rect 420 175 743 205
rect 392 169 743 175
rect 446 142 689 169
rect 473 115 689 142
<< ndiffc >>
rect 400 1265 420 1295
rect 370 1125 390 1155
<< pdiffc >>
rect 370 315 400 345
rect 400 175 420 205
<< psubdiff >>
rect 330 1375 410 1380
rect 330 1335 345 1375
rect 395 1335 410 1375
rect 330 1330 410 1335
<< nsubdiff >>
rect 335 135 405 140
rect 335 100 350 135
rect 390 100 405 135
rect 335 95 405 100
<< psubdiffcont >>
rect 345 1335 395 1375
<< nsubdiffcont >>
rect 350 100 390 135
<< polysilicon >>
rect 250 1181 365 1221
rect 770 1181 900 1221
rect 850 975 900 1181
rect 850 925 860 975
rect 890 925 900 975
rect 850 535 900 925
rect 850 485 860 535
rect 890 485 900 535
rect 850 295 900 485
rect 250 255 365 295
rect 770 255 900 295
<< polycontact >>
rect 860 925 890 975
rect 860 485 890 535
<< metal1 >>
rect 0 1400 1070 1440
rect 250 1240 290 1400
rect 330 1375 410 1380
rect 330 1335 345 1375
rect 395 1335 410 1375
rect 330 1305 410 1335
rect 310 1295 430 1305
rect 310 1270 320 1295
rect 345 1270 400 1295
rect 310 1265 400 1270
rect 420 1265 430 1295
rect 310 1255 430 1265
rect 250 1155 400 1165
rect 250 1125 370 1155
rect 390 1125 400 1155
rect 250 1115 400 1125
rect 250 355 300 1115
rect 850 975 900 995
rect 850 925 860 975
rect 890 925 900 975
rect 850 535 900 925
rect 850 485 860 535
rect 890 485 900 535
rect 850 455 900 485
rect 250 345 410 355
rect 250 315 370 345
rect 400 315 410 345
rect 250 305 410 315
rect 260 40 304 240
rect 340 205 430 215
rect 340 195 400 205
rect 340 175 345 195
rect 370 175 400 195
rect 420 175 430 205
rect 340 165 430 175
rect 335 135 405 165
rect 335 100 350 135
rect 390 100 405 135
rect 335 95 405 100
rect 0 0 1070 40
<< metal2 >>
rect 473 1330 689 1357
rect 446 1303 689 1330
rect 392 1249 743 1303
rect 365 1141 770 1249
rect 365 1114 446 1141
rect 365 1087 419 1114
rect 392 1060 419 1087
rect 527 1060 608 1141
rect 689 1114 770 1141
rect 716 1087 770 1114
rect 716 1060 743 1087
rect 392 1033 446 1060
rect 500 1033 635 1060
rect 689 1033 743 1060
rect 392 1006 554 1033
rect 581 1006 716 1033
rect 446 979 527 1006
rect 608 979 716 1006
rect 473 925 662 979
rect 311 898 392 925
rect 473 898 500 925
rect 527 898 554 925
rect 581 898 608 925
rect 635 898 662 925
rect 743 898 824 925
rect 284 844 419 898
rect 716 844 851 898
rect 311 817 473 844
rect 662 817 824 844
rect 392 790 500 817
rect 635 790 743 817
rect 446 763 554 790
rect 581 763 689 790
rect 500 709 635 763
rect 446 682 554 709
rect 581 682 689 709
rect 311 655 500 682
rect 635 655 851 682
rect 284 628 446 655
rect 689 628 851 655
rect 284 601 392 628
rect 743 601 851 628
rect 284 574 365 601
rect 770 574 851 601
rect 311 547 338 574
rect 473 547 500 574
rect 527 547 554 574
rect 581 547 608 574
rect 635 547 662 574
rect 797 547 824 574
rect 473 493 662 547
rect 446 466 527 493
rect 608 466 716 493
rect 392 439 554 466
rect 581 439 716 466
rect 392 412 446 439
rect 500 412 635 439
rect 689 412 743 439
rect 392 385 419 412
rect 365 358 419 385
rect 365 331 446 358
rect 527 331 608 412
rect 716 385 743 412
rect 716 358 770 385
rect 689 331 770 358
rect 365 223 770 331
rect 392 169 743 223
rect 446 142 689 169
rect 473 115 689 142
<< fillblock >>
rect 260 80 880 1390
<< labels >>
flabel metal1 s 250 1260 290 1305 0 FreeSans 240 90 0 0 VSS
port 1 nsew ground bidirectional abutment
flabel metal1 s 250 165 300 205 0 FreeSans 240 90 0 0 VDD
port 2 nsew power bidirectional abutment
flabel metal1 s 250 705 300 785 0 FreeSans 340 0 0 0 Y
port 3 s signal output
flabel metal1 s 850 705 900 785 0 FreeSans 340 0 0 0 A
port 4 e signal input
<< end >>
