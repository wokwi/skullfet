magic
tech gf180mcuC
magscale 1 2
timestamp 1670241224
<< metal1 >>
rect 14060 32300 18380 32840
rect 13520 31760 18380 32300
rect 12440 30680 19460 31760
rect 11900 28520 20000 30680
rect 11900 27980 13520 28520
rect 11900 27440 12980 27980
rect 12440 26900 12980 27440
rect 15140 26900 16760 28520
rect 18380 27980 20000 28520
rect 18920 27440 20000 27980
rect 18920 26900 19460 27440
rect 12440 26360 13520 26900
rect 14600 26360 17300 26900
rect 18380 26360 19460 26900
rect 12440 25820 15680 26360
rect 16220 25820 18920 26360
rect 13520 25280 15140 25820
rect 16760 25280 18920 25820
rect 14060 24200 17840 25280
rect 10820 23660 12440 24200
rect 14060 23660 14600 24200
rect 15140 23660 15680 24200
rect 16220 23660 16760 24200
rect 17300 23660 17840 24200
rect 19460 23660 21080 24200
rect 10280 22580 12980 23660
rect 18920 22580 21620 23660
rect 10820 22040 14060 22580
rect 17840 22040 21080 22580
rect 12440 21500 14600 22040
rect 17300 21500 19460 22040
rect 13520 20960 15680 21500
rect 16220 20960 18380 21500
rect 14600 19880 17300 20960
rect 13520 19340 15680 19880
rect 16220 19340 18380 19880
rect 10820 18800 14600 19340
rect 17300 18800 21620 19340
rect 10280 18260 13520 18800
rect 18380 18260 21620 18800
rect 10280 17720 12440 18260
rect 19460 17720 21620 18260
rect 10280 17180 11900 17720
rect 20000 17180 21620 17720
rect 10820 16640 11360 17180
rect 14060 16640 14600 17180
rect 15140 16640 15680 17180
rect 16220 16640 16760 17180
rect 17300 16640 17840 17180
rect 20540 16640 21080 17180
rect 14060 15560 17840 16640
rect 13520 15020 15140 15560
rect 16760 15020 18920 15560
rect 12440 14480 15680 15020
rect 16220 14480 18920 15020
rect 12440 13940 13520 14480
rect 14600 13940 17300 14480
rect 18380 13940 19460 14480
rect 12440 13400 12980 13940
rect 11900 12860 12980 13400
rect 11900 12320 13520 12860
rect 15140 12320 16760 13940
rect 18920 13400 19460 13940
rect 18920 12860 20000 13400
rect 18380 12320 20000 12860
rect 11900 10160 20000 12320
rect 12440 9080 19460 10160
rect 13520 8540 18380 9080
rect 14060 8000 18380 8540
rect 6800 6200 8400 6400
rect 9400 6200 9600 6400
rect 6600 6000 8400 6200
rect 9200 6000 9600 6200
rect 6400 4800 7000 6000
rect 7800 5600 8400 6000
rect 7800 5400 8200 5600
rect 7800 5200 8000 5400
rect 9000 5200 9600 6000
rect 10400 6200 10600 6400
rect 10200 6000 10800 6200
rect 10000 5800 10800 6000
rect 9800 5600 10600 5800
rect 9800 5400 10400 5600
rect 9800 5200 10200 5400
rect 9000 5000 10200 5200
rect 8800 4800 10000 5000
rect 6000 4600 8400 4800
rect 8600 4600 10000 4800
rect 6200 4400 8400 4600
rect 6800 3800 7000 4000
rect 6600 3600 7000 3800
rect 7800 3600 8400 4400
rect 9000 4400 10200 4600
rect 6400 3400 8200 3600
rect 6200 3200 8000 3400
rect 9000 3200 9600 4400
rect 9800 4200 10200 4400
rect 9800 4000 10400 4200
rect 9800 3800 10600 4000
rect 10000 3600 10800 3800
rect 10200 3400 10800 3600
rect 11000 3600 11600 6400
rect 12400 6200 12600 6400
rect 13600 6200 13800 6400
rect 15600 6200 15800 6400
rect 18000 6200 19600 6400
rect 20600 6200 22200 6400
rect 12400 6000 12800 6200
rect 13400 6000 13800 6200
rect 15400 6000 15800 6200
rect 17800 6000 19600 6200
rect 20400 6000 22200 6200
rect 23200 6000 23800 6400
rect 12400 3600 13000 6000
rect 13200 3600 13800 6000
rect 14800 3600 15000 3800
rect 11000 3400 12800 3600
rect 13200 3400 14200 3600
rect 14600 3400 15000 3600
rect 10400 3200 10600 3400
rect 11000 3200 12600 3400
rect 13200 3200 15000 3400
rect 15200 3600 15800 6000
rect 17600 5000 18200 6000
rect 19000 5600 19600 6000
rect 19000 5400 19400 5600
rect 19000 5200 19200 5400
rect 20200 5000 20800 6000
rect 21600 5600 22200 6000
rect 22400 5800 24400 6000
rect 22600 5600 24600 5800
rect 21600 5400 22000 5600
rect 23000 5400 24600 5600
rect 21600 5200 21800 5400
rect 17400 4800 18800 5000
rect 20000 4800 21400 5000
rect 17200 4600 18800 4800
rect 19800 4600 21400 4800
rect 16800 3600 17000 3800
rect 15200 3400 16200 3600
rect 16600 3400 17000 3600
rect 15200 3200 17000 3400
rect 17600 3200 18200 4600
rect 20200 3600 20800 4600
rect 21600 4200 21800 4400
rect 21600 4000 22000 4200
rect 21600 3600 22200 4000
rect 20200 3200 22200 3600
rect 23200 3600 23800 5400
rect 24200 5200 24600 5400
rect 24400 5000 24600 5200
rect 23200 3400 24200 3600
rect 23000 3200 24000 3400
rect 9000 3000 9200 3200
rect 13200 3000 13400 3200
rect 15200 3000 15400 3200
<< obsm2 >>
rect 10000 8000 22000 34000
rect 5000 2000 26000 8000
<< obsm3 >>
rect 10000 8000 22000 34000
rect 5000 2000 26000 8000
<< metal4 >>
rect 2000 2000 3000 34000
rect 14060 32300 18380 32840
rect 13520 31760 18380 32300
rect 12440 30680 19460 31760
rect 11900 28520 20000 30680
rect 11900 27980 13520 28520
rect 11900 27440 12980 27980
rect 12440 26900 12980 27440
rect 15140 26900 16760 28520
rect 18380 27980 20000 28520
rect 18920 27440 20000 27980
rect 18920 26900 19460 27440
rect 12440 26360 13520 26900
rect 14600 26360 17300 26900
rect 18380 26360 19460 26900
rect 12440 25820 15680 26360
rect 16220 25820 18920 26360
rect 13520 25280 15140 25820
rect 16760 25280 18920 25820
rect 14060 24200 17840 25280
rect 10820 23660 12440 24200
rect 14060 23660 14600 24200
rect 15140 23660 15680 24200
rect 16220 23660 16760 24200
rect 17300 23660 17840 24200
rect 19460 23660 21080 24200
rect 10280 22580 12980 23660
rect 18920 22580 21620 23660
rect 10820 22040 14060 22580
rect 17840 22040 21080 22580
rect 12440 21500 14600 22040
rect 17300 21500 19460 22040
rect 13520 20960 15680 21500
rect 16220 20960 18380 21500
rect 14600 19880 17300 20960
rect 13520 19340 15680 19880
rect 16220 19340 18380 19880
rect 10820 18800 14600 19340
rect 17300 18800 21620 19340
rect 10280 18260 13520 18800
rect 18380 18260 21620 18800
rect 10280 17720 12440 18260
rect 19460 17720 21620 18260
rect 10280 17180 11900 17720
rect 20000 17180 21620 17720
rect 10820 16640 11360 17180
rect 14060 16640 14600 17180
rect 15140 16640 15680 17180
rect 16220 16640 16760 17180
rect 17300 16640 17840 17180
rect 20540 16640 21080 17180
rect 14060 15560 17840 16640
rect 13520 15020 15140 15560
rect 16760 15020 18920 15560
rect 12440 14480 15680 15020
rect 16220 14480 18920 15020
rect 12440 13940 13520 14480
rect 14600 13940 17300 14480
rect 18380 13940 19460 14480
rect 12440 13400 12980 13940
rect 11900 12860 12980 13400
rect 11900 12320 13520 12860
rect 15140 12320 16760 13940
rect 18920 13400 19460 13940
rect 18920 12860 20000 13400
rect 18380 12320 20000 12860
rect 11900 10160 20000 12320
rect 12440 9080 19460 10160
rect 13520 8540 18380 9080
rect 14060 8000 18380 8540
rect 6800 6200 8400 6400
rect 9400 6200 9600 6400
rect 6600 6000 8400 6200
rect 9200 6000 9600 6200
rect 6400 4800 7000 6000
rect 7800 5600 8400 6000
rect 7800 5400 8200 5600
rect 7800 5200 8000 5400
rect 9000 5200 9600 6000
rect 10400 6200 10600 6400
rect 10200 6000 10800 6200
rect 10000 5800 10800 6000
rect 9800 5600 10600 5800
rect 9800 5400 10400 5600
rect 9800 5200 10200 5400
rect 9000 5000 10200 5200
rect 8800 4800 10000 5000
rect 6000 4600 8400 4800
rect 8600 4600 10000 4800
rect 6200 4400 8400 4600
rect 6800 3800 7000 4000
rect 6600 3600 7000 3800
rect 7800 3600 8400 4400
rect 9000 4400 10200 4600
rect 6400 3400 8200 3600
rect 6200 3200 8000 3400
rect 9000 3200 9600 4400
rect 9800 4200 10200 4400
rect 9800 4000 10400 4200
rect 9800 3800 10600 4000
rect 10000 3600 10800 3800
rect 10200 3400 10800 3600
rect 11000 3600 11600 6400
rect 12400 6200 12600 6400
rect 13600 6200 13800 6400
rect 15600 6200 15800 6400
rect 18000 6200 19600 6400
rect 20600 6200 22200 6400
rect 12400 6000 12800 6200
rect 13400 6000 13800 6200
rect 15400 6000 15800 6200
rect 17800 6000 19600 6200
rect 20400 6000 22200 6200
rect 23200 6000 23800 6400
rect 12400 3600 13000 6000
rect 13200 3600 13800 6000
rect 14800 3600 15000 3800
rect 11000 3400 12800 3600
rect 13200 3400 14200 3600
rect 14600 3400 15000 3600
rect 10400 3200 10600 3400
rect 11000 3200 12600 3400
rect 13200 3200 15000 3400
rect 15200 3600 15800 6000
rect 17600 5000 18200 6000
rect 19000 5600 19600 6000
rect 19000 5400 19400 5600
rect 19000 5200 19200 5400
rect 20200 5000 20800 6000
rect 21600 5600 22200 6000
rect 22400 5800 24400 6000
rect 22600 5600 24600 5800
rect 21600 5400 22000 5600
rect 23000 5400 24600 5600
rect 21600 5200 21800 5400
rect 17400 4800 18800 5000
rect 20000 4800 21400 5000
rect 17200 4600 18800 4800
rect 19800 4600 21400 4800
rect 16800 3600 17000 3800
rect 15200 3400 16200 3600
rect 16600 3400 17000 3600
rect 15200 3200 17000 3400
rect 17600 3200 18200 4600
rect 20200 3600 20800 4600
rect 21600 4200 21800 4400
rect 21600 4000 22000 4200
rect 21600 3600 22200 4000
rect 20200 3200 22200 3600
rect 23200 3600 23800 5400
rect 24200 5200 24600 5400
rect 24400 5000 24600 5200
rect 23200 3400 24200 3600
rect 23000 3200 24000 3400
rect 9000 3000 9200 3200
rect 13200 3000 13400 3200
rect 15200 3000 15400 3200
rect 29000 2000 30000 34000
<< labels >>
flabel metal4 s 29000 33000 30000 34000 0 FreeSans 240 0 0 0 vss
port 1 nsew ground bidirectional abutment
flabel metal4 s 2000 33000 3000 34000 0 FreeSans 240 0 0 0 vdd
port 2 nsew power bidirectional abutment
<< end >>
