magic
tech sky130A
timestamp 1640345212
<< nwell >>
rect 75 -1405 595 -835
<< pwell >>
rect 75 -590 595 -75
<< nmos >>
rect 135 -284 540 -244
<< pmos >>
rect 135 -1210 540 -1170
<< ndiff >>
rect 243 -135 459 -108
rect 216 -162 459 -135
rect 162 -170 513 -162
rect 162 -200 170 -170
rect 190 -200 513 -170
rect 162 -216 513 -200
rect 135 -244 540 -216
rect 135 -310 540 -284
rect 135 -340 140 -310
rect 160 -324 540 -310
rect 160 -340 216 -324
rect 135 -351 216 -340
rect 135 -378 189 -351
rect 162 -405 189 -378
rect 297 -405 378 -324
rect 459 -351 540 -324
rect 486 -378 540 -351
rect 486 -405 513 -378
rect 162 -432 216 -405
rect 270 -432 405 -405
rect 459 -432 513 -405
rect 162 -459 324 -432
rect 351 -459 486 -432
rect 216 -486 297 -459
rect 378 -486 486 -459
rect 243 -540 432 -486
rect 243 -567 270 -540
rect 297 -567 324 -540
rect 351 -567 378 -540
rect 405 -567 432 -540
<< pdiff >>
rect 243 -918 270 -891
rect 297 -918 324 -891
rect 351 -918 378 -891
rect 405 -918 432 -891
rect 243 -972 432 -918
rect 216 -999 297 -972
rect 378 -999 486 -972
rect 162 -1026 324 -999
rect 351 -1026 486 -999
rect 162 -1053 216 -1026
rect 270 -1053 405 -1026
rect 459 -1053 513 -1026
rect 162 -1080 189 -1053
rect 135 -1107 189 -1080
rect 135 -1120 216 -1107
rect 135 -1150 140 -1120
rect 170 -1134 216 -1120
rect 297 -1134 378 -1053
rect 486 -1080 513 -1053
rect 486 -1107 540 -1080
rect 459 -1134 540 -1107
rect 170 -1150 540 -1134
rect 135 -1170 540 -1150
rect 135 -1242 540 -1210
rect 162 -1260 513 -1242
rect 162 -1290 170 -1260
rect 190 -1290 513 -1260
rect 162 -1296 513 -1290
rect 216 -1323 459 -1296
rect 243 -1350 459 -1323
<< ndiffc >>
rect 170 -200 190 -170
rect 140 -340 160 -310
<< pdiffc >>
rect 140 -1150 170 -1120
rect 170 -1290 190 -1260
<< psubdiff >>
rect 100 -90 180 -85
rect 100 -130 115 -90
rect 165 -130 180 -90
rect 100 -135 180 -130
<< nsubdiff >>
rect 105 -1330 175 -1325
rect 105 -1365 120 -1330
rect 160 -1365 175 -1330
rect 105 -1370 175 -1365
<< psubdiffcont >>
rect 115 -130 165 -90
<< nsubdiffcont >>
rect 120 -1365 160 -1330
<< poly >>
rect 20 -284 135 -244
rect 540 -284 670 -244
rect 620 -490 670 -284
rect 620 -540 630 -490
rect 660 -540 670 -490
rect 620 -930 670 -540
rect 620 -980 630 -930
rect 660 -980 670 -930
rect 620 -1170 670 -980
rect 20 -1210 135 -1170
rect 540 -1210 670 -1170
<< polycont >>
rect 630 -540 660 -490
rect 630 -980 660 -930
<< locali >>
rect 100 -90 180 -85
rect 100 -130 115 -90
rect 165 -130 180 -90
rect 100 -160 180 -130
rect 80 -170 200 -160
rect 80 -200 90 -170
rect 120 -200 170 -170
rect 190 -200 200 -170
rect 80 -210 200 -200
rect 20 -310 170 -300
rect 20 -340 140 -310
rect 160 -340 170 -310
rect 20 -350 170 -340
rect 20 -1110 70 -350
rect 620 -490 670 -470
rect 620 -540 630 -490
rect 660 -540 670 -490
rect 620 -930 670 -540
rect 620 -980 630 -930
rect 660 -980 670 -930
rect 620 -1010 670 -980
rect 20 -1120 180 -1110
rect 20 -1150 140 -1120
rect 170 -1150 180 -1120
rect 20 -1160 180 -1150
rect 110 -1260 200 -1250
rect 110 -1290 120 -1260
rect 150 -1290 170 -1260
rect 190 -1290 200 -1260
rect 110 -1300 200 -1290
rect 105 -1330 175 -1300
rect 105 -1365 120 -1330
rect 160 -1365 175 -1330
rect 105 -1370 175 -1365
<< viali >>
rect 90 -200 120 -170
rect 120 -1290 150 -1260
<< metal1 >>
rect 20 -170 130 -160
rect 20 -200 90 -170
rect 120 -200 130 -170
rect 20 -210 130 -200
rect 81 -567 162 -540
rect 513 -567 594 -540
rect 54 -621 189 -567
rect 486 -621 621 -567
rect 81 -648 243 -621
rect 432 -648 594 -621
rect 162 -675 270 -648
rect 405 -675 513 -648
rect 216 -702 324 -675
rect 351 -702 459 -675
rect 270 -756 405 -702
rect 216 -783 324 -756
rect 351 -783 459 -756
rect 81 -810 270 -783
rect 405 -810 621 -783
rect 54 -837 216 -810
rect 459 -837 621 -810
rect 54 -864 162 -837
rect 513 -864 621 -837
rect 54 -891 135 -864
rect 540 -891 621 -864
rect 81 -918 108 -891
rect 567 -918 594 -891
rect 20 -1260 160 -1250
rect 20 -1290 120 -1260
rect 150 -1290 160 -1260
rect 20 -1300 160 -1290
<< labels >>
flabel metal1 s 20 -210 70 -160 0 FreeSans 240 90 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 20 -1300 70 -1250 0 FreeSans 240 90 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 20 -760 70 -680 0 FreeSans 340 0 0 0 Y
port 3 s signal output
flabel locali s 620 -760 670 -680 0 FreeSans 340 0 0 0 A
port 4 e signal input
flabel metal1 s 80 -1300 130 -1250 0 FreeSans 240 90 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 80 -210 130 -160 0 FreeSans 240 90 0 0 VNB
port 6 nsew ground bidirectional
<< end >>
