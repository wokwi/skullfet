magic
tech sky130A
magscale 1 2
timestamp 1640713472
<< nwell >>
rect 1242 -1728 2295 -972
rect 189 -1944 2295 -1728
rect 189 -2781 1161 -1944
<< nmos >>
rect 270 -594 1080 -486
rect -594 -1836 -486 -1026
<< pmos >>
rect 1836 -1836 1944 -1026
rect 270 -2430 1080 -2322
<< ndiff >>
rect 486 -270 918 -216
rect 432 -324 918 -270
rect 324 -351 1026 -324
rect 324 -405 351 -351
rect 405 -405 1026 -351
rect 324 -432 1026 -405
rect 270 -486 1080 -432
rect 270 -648 1080 -594
rect 270 -702 432 -648
rect 270 -756 378 -702
rect 324 -810 378 -756
rect 594 -810 756 -648
rect 918 -702 999 -648
rect 1053 -702 1080 -648
rect 972 -756 1080 -702
rect 972 -810 1026 -756
rect 324 -864 432 -810
rect 540 -864 810 -810
rect 918 -864 1026 -810
rect 324 -918 648 -864
rect 702 -918 972 -864
rect 432 -972 594 -918
rect 756 -972 972 -918
rect -648 -1080 -594 -1026
rect -756 -1188 -594 -1080
rect -864 -1620 -594 -1188
rect -810 -1674 -594 -1620
rect -756 -1701 -594 -1674
rect -756 -1755 -729 -1701
rect -675 -1755 -594 -1701
rect -756 -1782 -594 -1755
rect -648 -1836 -594 -1782
rect -486 -1053 -324 -1026
rect -486 -1107 -432 -1053
rect -378 -1080 -324 -1053
rect 486 -1080 864 -972
rect -378 -1107 -216 -1080
rect -486 -1134 -216 -1107
rect 486 -1134 540 -1080
rect 594 -1134 648 -1080
rect 702 -1134 756 -1080
rect 810 -1134 864 -1080
rect -486 -1188 -378 -1134
rect -270 -1188 -108 -1134
rect -486 -1350 -432 -1188
rect -216 -1242 -108 -1188
rect -216 -1296 54 -1242
rect -270 -1350 0 -1296
rect -486 -1404 -162 -1350
rect -108 -1404 54 -1350
rect -486 -1458 -216 -1404
rect -108 -1458 0 -1404
rect -486 -1512 -162 -1458
rect -108 -1512 54 -1458
rect -486 -1674 -432 -1512
rect -270 -1566 0 -1512
rect -216 -1620 54 -1566
rect -216 -1674 -108 -1620
rect -486 -1728 -378 -1674
rect -270 -1728 -162 -1674
rect -486 -1782 -162 -1728
rect -486 -1836 -324 -1782
<< pdiff >>
rect 1674 -1053 1836 -1026
rect 1674 -1080 1728 -1053
rect 1512 -1107 1728 -1080
rect 1782 -1107 1836 -1053
rect 1512 -1134 1836 -1107
rect 1512 -1188 1620 -1134
rect 1728 -1188 1836 -1134
rect 1458 -1242 1566 -1188
rect 1296 -1296 1566 -1242
rect 1350 -1350 1620 -1296
rect 1782 -1350 1836 -1188
rect 1296 -1404 1458 -1350
rect 1512 -1404 1836 -1350
rect 1350 -1458 1458 -1404
rect 1566 -1458 1836 -1404
rect 1296 -1512 1458 -1458
rect 1512 -1512 1836 -1458
rect 1350 -1566 1620 -1512
rect 1296 -1620 1566 -1566
rect 1458 -1674 1566 -1620
rect 1782 -1674 1836 -1512
rect 1458 -1728 1620 -1674
rect 1728 -1728 1836 -1674
rect 1566 -1755 1836 -1728
rect 1566 -1782 1728 -1755
rect 486 -1836 540 -1782
rect 594 -1836 648 -1782
rect 702 -1836 756 -1782
rect 810 -1836 864 -1782
rect 1674 -1809 1728 -1782
rect 1782 -1809 1836 -1755
rect 1674 -1836 1836 -1809
rect 1944 -1080 1998 -1026
rect 1944 -1188 2106 -1080
rect 1944 -1242 2160 -1188
rect 1944 -1674 2214 -1242
rect 1944 -1701 2106 -1674
rect 1944 -1755 2025 -1701
rect 2079 -1755 2106 -1701
rect 1944 -1782 2106 -1755
rect 1944 -1836 1998 -1782
rect 486 -1944 864 -1836
rect 432 -1998 594 -1944
rect 756 -1998 972 -1944
rect 324 -2052 648 -1998
rect 702 -2052 972 -1998
rect 324 -2106 432 -2052
rect 540 -2106 810 -2052
rect 918 -2106 1026 -2052
rect 324 -2160 378 -2106
rect 270 -2214 378 -2160
rect 270 -2268 432 -2214
rect 594 -2268 756 -2106
rect 972 -2160 1026 -2106
rect 972 -2214 1080 -2160
rect 918 -2268 999 -2214
rect 1053 -2268 1080 -2214
rect 270 -2322 1080 -2268
rect 270 -2484 1080 -2430
rect 324 -2511 1026 -2484
rect 324 -2565 945 -2511
rect 999 -2565 1026 -2511
rect 324 -2592 1026 -2565
rect 432 -2646 918 -2592
rect 486 -2700 918 -2646
<< ndiffc >>
rect 351 -405 405 -351
rect 999 -702 1053 -648
rect -729 -1755 -675 -1701
rect -432 -1107 -378 -1053
<< pdiffc >>
rect 1728 -1107 1782 -1053
rect 1728 -1809 1782 -1755
rect 2025 -1755 2079 -1701
rect 999 -2268 1053 -2214
rect 945 -2565 999 -2511
<< psubdiff >>
rect -918 -1755 -810 -1728
rect -918 -1836 -864 -1755
rect -918 -1863 -810 -1836
<< nsubdiff >>
rect 2160 -1755 2241 -1728
rect 2214 -1836 2241 -1755
rect 2160 -1890 2241 -1836
rect 972 -2700 999 -2646
rect 1080 -2700 1107 -2646
rect 972 -2727 1107 -2700
<< psubdiffcont >>
rect -864 -1836 -810 -1755
<< nsubdiffcont >>
rect 2160 -1836 2214 -1755
rect 999 -2700 1080 -2646
<< poly >>
rect 108 -594 270 -486
rect 1080 -513 1944 -486
rect 1080 -567 1431 -513
rect 1485 -567 1863 -513
rect 1917 -567 1944 -513
rect 1080 -594 1944 -567
rect -594 -1026 -486 -864
rect 1836 -1026 1944 -594
rect -594 -2322 -486 -1836
rect 1836 -1998 1944 -1836
rect -594 -2349 270 -2322
rect -594 -2403 -567 -2349
rect -513 -2403 -135 -2349
rect -81 -2403 270 -2349
rect -594 -2430 270 -2403
rect 1080 -2430 1242 -2322
<< polycont >>
rect 1431 -567 1485 -513
rect 1863 -567 1917 -513
rect -567 -2403 -513 -2349
rect -135 -2403 -81 -2349
<< locali >>
rect -459 -351 405 -324
rect -459 -405 351 -351
rect -459 -432 405 -405
rect -459 -1053 -351 -432
rect 1404 -513 1944 -486
rect 1404 -567 1431 -513
rect 1485 -567 1863 -513
rect 1917 -567 1944 -513
rect 1404 -594 1944 -567
rect 999 -648 1350 -621
rect 1053 -702 1350 -648
rect 999 -729 1350 -702
rect 1242 -837 1809 -729
rect -459 -1107 -432 -1053
rect -378 -1107 -351 -1053
rect 1701 -1053 1809 -837
rect 1701 -1107 1728 -1053
rect 1782 -1107 1809 -1053
rect -864 -1755 -729 -1701
rect -675 -1755 -648 -1701
rect 1998 -1755 2025 -1701
rect 2079 -1728 2106 -1701
rect 2079 -1755 2214 -1728
rect -810 -1836 -648 -1755
rect -864 -1863 -648 -1836
rect -756 -2484 -648 -1863
rect 1701 -1809 1728 -1755
rect 1782 -1809 1809 -1755
rect 1701 -2187 1809 -1809
rect 999 -2214 1809 -2187
rect 1053 -2268 1809 -2214
rect 999 -2295 1809 -2268
rect 1998 -1836 2160 -1755
rect 1998 -1863 2214 -1836
rect -594 -2349 -54 -2322
rect -594 -2403 -567 -2349
rect -513 -2403 -135 -2349
rect -81 -2403 -54 -2349
rect -594 -2430 -54 -2403
rect 1998 -2403 2106 -1863
rect -756 -2592 -729 -2484
rect 945 -2511 1404 -2484
rect 999 -2565 1404 -2511
rect 945 -2592 1404 -2565
rect 1485 -2592 2106 -2484
rect 945 -2646 1134 -2592
rect 945 -2700 999 -2646
rect 1080 -2700 1134 -2646
<< viali >>
rect 1998 -2484 2106 -2403
rect -729 -2592 -648 -2484
rect 1404 -2592 1485 -2484
<< metal1 >>
rect 486 -270 918 -216
rect 432 -324 918 -270
rect 324 -432 1026 -324
rect 270 -648 1080 -432
rect 270 -702 432 -648
rect 270 -756 378 -702
rect 324 -810 378 -756
rect 594 -810 756 -648
rect 918 -702 1080 -648
rect 972 -756 1080 -702
rect 972 -810 1026 -756
rect 324 -864 432 -810
rect 540 -864 810 -810
rect 918 -864 1026 -810
rect 324 -918 648 -864
rect 702 -918 972 -864
rect 432 -972 594 -918
rect 756 -972 972 -918
rect -648 -1080 -324 -1026
rect 486 -1080 864 -972
rect 1674 -1080 1998 -1026
rect -756 -1134 -216 -1080
rect 162 -1134 324 -1080
rect 486 -1134 540 -1080
rect 594 -1134 648 -1080
rect 702 -1134 756 -1080
rect 810 -1134 864 -1080
rect 1026 -1134 1188 -1080
rect 1512 -1134 2106 -1080
rect -756 -1188 -378 -1134
rect -270 -1188 -108 -1134
rect -864 -1350 -432 -1188
rect -216 -1242 -108 -1188
rect 108 -1242 378 -1134
rect 972 -1242 1242 -1134
rect 1512 -1188 1620 -1134
rect 1728 -1188 2106 -1134
rect 1458 -1242 1566 -1188
rect -216 -1296 54 -1242
rect 162 -1296 486 -1242
rect 864 -1296 1188 -1242
rect 1296 -1296 1566 -1242
rect 1782 -1242 2160 -1188
rect -270 -1350 0 -1296
rect 324 -1350 540 -1296
rect 810 -1350 1026 -1296
rect 1350 -1350 1620 -1296
rect 1782 -1350 2214 -1242
rect -864 -1404 -162 -1350
rect -108 -1404 54 -1350
rect 432 -1404 648 -1350
rect 702 -1404 918 -1350
rect 1296 -1404 1458 -1350
rect 1512 -1404 2214 -1350
rect -864 -1458 -216 -1404
rect -108 -1458 0 -1404
rect -864 -1512 -162 -1458
rect -108 -1512 54 -1458
rect 540 -1512 810 -1404
rect 1350 -1458 1458 -1404
rect 1566 -1458 2214 -1404
rect 1296 -1512 1458 -1458
rect 1512 -1512 2214 -1458
rect -864 -1620 -432 -1512
rect -270 -1566 0 -1512
rect 432 -1566 648 -1512
rect 702 -1566 918 -1512
rect 1350 -1566 1620 -1512
rect -810 -1674 -432 -1620
rect -216 -1620 54 -1566
rect 162 -1620 540 -1566
rect 810 -1620 1242 -1566
rect 1296 -1620 1566 -1566
rect -216 -1674 -108 -1620
rect 108 -1674 432 -1620
rect 918 -1674 1242 -1620
rect -756 -1728 -378 -1674
rect -270 -1728 -162 -1674
rect -756 -1782 -162 -1728
rect 108 -1728 324 -1674
rect 1026 -1728 1242 -1674
rect 1458 -1674 1566 -1620
rect 1782 -1674 2214 -1512
rect 1458 -1728 1620 -1674
rect 1728 -1728 2106 -1674
rect 108 -1782 270 -1728
rect 1080 -1782 1242 -1728
rect 1566 -1782 2106 -1728
rect -648 -1836 -324 -1782
rect 162 -1836 216 -1782
rect 486 -1836 540 -1782
rect 594 -1836 648 -1782
rect 702 -1836 756 -1782
rect 810 -1836 864 -1782
rect 1134 -1836 1188 -1782
rect 1674 -1836 1998 -1782
rect 486 -1944 864 -1836
rect 432 -1998 594 -1944
rect 756 -1998 972 -1944
rect 324 -2052 648 -1998
rect 702 -2052 972 -1998
rect 324 -2106 432 -2052
rect 540 -2106 810 -2052
rect 918 -2106 1026 -2052
rect 324 -2160 378 -2106
rect 270 -2214 378 -2160
rect 270 -2268 432 -2214
rect 594 -2268 756 -2106
rect 972 -2160 1026 -2106
rect 972 -2214 1080 -2160
rect 918 -2268 1080 -2214
rect -756 -2484 -324 -2457
rect 270 -2484 1080 -2268
rect 1377 -2403 2187 -2376
rect 1377 -2484 1998 -2403
rect 2106 -2484 2187 -2403
rect -756 -2592 -729 -2484
rect -648 -2592 -324 -2484
rect 324 -2592 1026 -2484
rect 1377 -2592 1404 -2484
rect 1485 -2592 2187 -2484
rect -756 -2619 -324 -2592
rect -756 -2781 -648 -2619
rect 432 -2646 918 -2592
rect 1377 -2646 2187 -2592
rect 486 -2700 918 -2646
rect -945 -2862 1998 -2781
rect 2079 -2916 2187 -2646
rect -945 -2997 2187 -2916
<< metal2 >>
rect 486 -270 918 -216
rect 432 -324 918 -270
rect 324 -432 1026 -324
rect 270 -648 1080 -432
rect 270 -702 432 -648
rect 270 -756 378 -702
rect 324 -810 378 -756
rect 594 -810 756 -648
rect 918 -702 1080 -648
rect 972 -756 1080 -702
rect 972 -810 1026 -756
rect 324 -864 432 -810
rect 540 -864 810 -810
rect 918 -864 1026 -810
rect 324 -918 648 -864
rect 702 -918 972 -864
rect 432 -972 594 -918
rect 756 -972 972 -918
rect -648 -1080 -324 -1026
rect 486 -1080 864 -972
rect 1674 -1080 1998 -1026
rect -756 -1134 -216 -1080
rect 486 -1134 540 -1080
rect 594 -1134 648 -1080
rect 702 -1134 756 -1080
rect 810 -1134 864 -1080
rect 1512 -1134 2106 -1080
rect -756 -1188 -378 -1134
rect -270 -1188 -108 -1134
rect 1512 -1188 1620 -1134
rect 1728 -1188 2106 -1134
rect -864 -1350 -432 -1188
rect -216 -1242 -108 -1188
rect 1458 -1242 1566 -1188
rect -216 -1296 54 -1242
rect 1296 -1296 1566 -1242
rect 1782 -1242 2160 -1188
rect -270 -1350 0 -1296
rect 1350 -1350 1620 -1296
rect 1782 -1350 2214 -1242
rect -864 -1404 -162 -1350
rect -108 -1404 54 -1350
rect 1296 -1404 1458 -1350
rect 1512 -1404 2214 -1350
rect -864 -1458 -216 -1404
rect -108 -1458 0 -1404
rect 1350 -1458 1458 -1404
rect 1566 -1458 2214 -1404
rect -864 -1512 -162 -1458
rect -108 -1512 54 -1458
rect 1296 -1512 1458 -1458
rect 1512 -1512 2214 -1458
rect -864 -1620 -432 -1512
rect -270 -1566 0 -1512
rect 1350 -1566 1620 -1512
rect -810 -1674 -432 -1620
rect -216 -1620 54 -1566
rect 1296 -1620 1566 -1566
rect -216 -1674 -108 -1620
rect 1458 -1674 1566 -1620
rect 1782 -1674 2214 -1512
rect -756 -1728 -378 -1674
rect -270 -1728 -162 -1674
rect 1458 -1728 1620 -1674
rect 1728 -1728 2106 -1674
rect -756 -1782 -162 -1728
rect 1566 -1782 2106 -1728
rect -648 -1836 -324 -1782
rect 486 -1836 540 -1782
rect 594 -1836 648 -1782
rect 702 -1836 756 -1782
rect 810 -1836 864 -1782
rect 1674 -1836 1998 -1782
rect 486 -1944 864 -1836
rect 432 -1998 594 -1944
rect 756 -1998 972 -1944
rect 324 -2052 648 -1998
rect 702 -2052 972 -1998
rect 324 -2106 432 -2052
rect 540 -2106 810 -2052
rect 918 -2106 1026 -2052
rect 324 -2160 378 -2106
rect 270 -2214 378 -2160
rect 270 -2268 432 -2214
rect 594 -2268 756 -2106
rect 972 -2160 1026 -2106
rect 972 -2214 1080 -2160
rect 918 -2268 1080 -2214
rect 270 -2484 1080 -2268
rect 324 -2592 1026 -2484
rect 432 -2646 918 -2592
rect 486 -2700 918 -2646
<< labels >>
flabel locali s 1566 -594 1755 -486 0 FreeSans 240 0 0 0 A
port 1 nsew signal input
flabel locali s -405 -2430 -216 -2322 0 FreeSans 240 0 0 0 B
port 2 nsew signal input
flabel locali s 1431 -837 1620 -729 0 FreeSans 240 0 0 0 Y
port 3 nsew signal output
flabel metal1 s 1701 -2592 1890 -2484 0 FreeSans 240 0 0 0 VPWR
port 4 nsew power bidirectional
flabel metal1 s -756 -2781 -648 -2619 0 FreeSans 240 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1242 -2592 1350 -2484 0 FreeSans 240 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s -756 -2187 -648 -2079 0 FreeSans 240 0 0 0 VNB
port 7 nsew ground bidirectional
<< end >>
